* FILE: project.sp

********************** begin header *****************************

* Sample Spice Header file for Generic 2.5V 0.25 um process (mmi25)

.OPTIONS post NOMOD post_version=9601

**################################################
* Only Typical/Typical spice models included
.include '${MMI_TOOLS}/sue/schematics/mspice/mmi25.mod'
* NOTE: these are contrived spice models
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=0,2,10,12 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3,13 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.6u
.param lp_min   =  0.6u

* used in source/drain area/perimeter calculation
.param sdd        =  0.66

.PARAM vddp=2.25	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "project" generated by MMI_SUE5.6.18 on Wed Dec 02 
*+ 11:44:58 CST 2015.

.SUBCKT nand A B Y 
M_1 net_1 A gnd gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' 
+ as='arean(1,sdd)' pd='perin(1,sdd)' ps='perin(1,sdd)' 
M_2 Y B net_1 gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' 
+ as='arean(1,sdd)' pd='perin(1,sdd)' ps='perin(1,sdd)' 
M_3 Y A vdd vdd p W='2*1u' L=lp_min ad='areap(2,sdd)' as='areap(2,sdd)' 
+ pd='perip(2,sdd)' ps='perip(2,sdd)' 
M_4 Y B vdd vdd p W='2*1u' L=lp_min ad='areap(2,sdd)' as='areap(2,sdd)' 
+ pd='perip(2,sdd)' ps='perip(2,sdd)' 
.ENDS	$ nand

.SUBCKT inv A Y 
M_1 Y A gnd gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' as='arean(1,sdd)' 
+ pd='perin(1,sdd)' ps='perin(1,sdd)' 
M_2 Y A vdd vdd p W='2*1u' L=lp_min ad='areap(2,sdd)' as='areap(2,sdd)' 
+ pd='perip(2,sdd)' ps='perip(2,sdd)' 
.ENDS	$ inv

.SUBCKT inverter in out WP=2 LP=lp_min WN=1 LN=ln_min
M_1 out in gnd gnd n W='WN*1u' L=LN ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_2 out in vdd vdd p W='WP*1u' L=LP ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
.ENDS	$ inverter

.SUBCKT nand2 in0 in1 out WP=2 WN=2
M_1 out in0 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_2 out in0 net_1 gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_3 out in1 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_4 net_1 in1 gnd gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
.ENDS	$ nand2

.SUBCKT 21mux A B Out S 
Xnand2 B S net_1 nand2 
Xnand2_1 net_3 A net_2 nand2 
Xnand2_2 net_1 net_2 Out nand2 
Xinverter S net_3 inverter 
.ENDS	$ 21mux

.SUBCKT dffpos Clk D Q 
M_1 net_10 net_1 gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_2 net_4 Clk net_10 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_3 net_1 net_4 gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_4 net_4 Clk_b net_6 vdd p W='3*1u' L=lp_min ad='areap(3,sdd)' 
+ as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_5 net_6 net_1 vdd vdd p W='3*1u' L=lp_min ad='areap(3,sdd)' 
+ as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_6 Clk_b Clk gnd gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_7 Clk_b Clk vdd vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_8 net_5 net_1 gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_9 net_3 Clk net_5 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_10 net_3 Clk_b net_9 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_11 net_9 net_1 vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_12 net_1 net_4 vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_13 Q net_3 gnd gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_14 Q net_3 vdd vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_15 net_2 D gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_16 net_4 Clk_b net_2 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_17 net_4 Clk net_8 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_18 net_8 D vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_19 net_11 Q gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_20 net_3 Clk_b net_11 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_21 net_3 Clk net_7 vdd p W='3*1u' L=lp_min ad='areap(3,sdd)' 
+ as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_22 net_7 Q vdd vdd p W='3*1u' L=lp_min ad='areap(3,sdd)' 
+ as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
.ENDS	$ dffpos

.SUBCKT FA a b c cout sum 
M_1 net_10 net_2 net_9 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_2 net_9 a gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_3 net_9 b gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_4 net_9 c gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_5 net_10 c net_12 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_6 net_12 b net_8 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_7 net_8 a gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_8 net_2 c net_5 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_9 net_5 a gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_10 net_5 b gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_11 net_2 b net_4 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_12 net_4 a gnd gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_13 net_11 a vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_14 net_11 b vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_15 net_11 c vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_16 net_10 net_2 net_11 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_17 net_1 b net_3 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_18 net_10 c net_1 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_19 net_3 a vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_20 net_6 a vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_21 net_6 b vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_22 net_2 c net_6 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_23 net_2 b net_7 vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
M_24 net_7 a vdd vdd p W='6*1u' L=lp_min ad='areap(6,sdd)' 
+ as='areap(6,sdd)' pd='perip(6,sdd)' ps='perip(6,sdd)' 
Xinv net_2 cout inv 
Xinv_1 net_10 sum inv 
.ENDS	$ FA

.SUBCKT xor2 a b out 
M_1 net_4 b vdd vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_2 out net_1 net_4 vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_3 out a net_6 vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_4 net_6 net_3 vdd vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_5 net_2 b gnd gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_6 net_5 net_3 gnd gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_7 out a net_2 gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_8 out net_1 net_5 gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_9 net_1 a vdd vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_10 net_1 a gnd gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
M_11 net_3 b vdd vdd p W='12*1u' L=lp_min ad='areap(12,sdd)' 
+ as='areap(12,sdd)' pd='perip(12,sdd)' ps='perip(12,sdd)' 
M_12 net_3 b gnd gnd n W='6*1u' L=ln_min ad='arean(6,sdd)' 
+ as='arean(6,sdd)' pd='perin(6,sdd)' ps='perin(6,sdd)' 
.ENDS	$ xor2

.SUBCKT bitslice A B Cin Clk Cout Out S subtract 
Xxor2 A subtract net_2 xor2 
X21mux Out B net_1 S 21mux 
XFA net_2 net_1 Cin Cout net_3 FA 
Xdffpos Clk net_3 Out dffpos 
.ENDS	$ bitslice

* start main CELL project
* .SUBCKT project A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] B[0] B[1] B[2] 
*+ B[3] B[4] B[5] B[6] B[7] Clk Cout Out[0] Out[1] Out[2] Out[3] Out[4] 
*+ Out[5] Out[6] Out[7] S loadR subtract 
Xnand loadR Clk net_9 nand 
Xinv net_9 net_1 inv 
Xbitslice A[3] B[3] net_3 net_1 net_2 Out[3] S subtract bitslice 
Xbitslice_1 A[4] B[4] net_2 net_1 net_5 uc_net_10 S subtract bitslice 
Xbitslice_2 A[5] B[5] net_5 net_1 net_6 Out[5] S subtract bitslice 
Xbitslice_3 A[2] B[2] net_4 net_1 net_3 Out[2] S subtract bitslice 
Xbitslice_4 A[6] B[6] net_6 net_1 net_7 Out[6] S subtract bitslice 
Xbitslice_5 A[7] B[7] net_7 net_1 Cout Out[7] S subtract bitslice 
Xbitslice_6 A[1] B[1] net_8 net_1 net_4 Out[1] S subtract bitslice 
Xbitslice_7 A[0] B[0] subtract net_1 net_8 Out[0] S subtract bitslice 
* .ENDS	$ project

.GLOBAL gnd vdd

.END

