* SPICE3 file created from mux21.ext - technology: scmos

.option scale=0.3u

M1000 nand_1/A A nand_2/vdd nand_2/vdd pfet w=20 l=2
+  ad=120 pd=52 as=300 ps=150
M1001 nand_2/vdd S' nand_1/A nand_2/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 nand_2/a_9_6# A nand_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=350 ps=180
M1003 nand_1/A S' nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 S' nand_0/A nand_2/vdd nand_2/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1005 S' nand_0/A nand_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1006 out nand_1/A nand_0/vdd nand_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=400 ps=200
M1007 nand_0/vdd nand_1/B out nand_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 nand_1/a_9_6# nand_1/A nand_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1009 out nand_1/B nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1010 nand_1/B nand_0/A nand_0/vdd nand_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1011 nand_0/vdd B nand_1/B nand_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 nand_0/a_9_6# nand_0/A nand_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1013 nand_1/B B nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 S' nand_2/vdd 5.711850fF
C1 nand_0/vdd nand_1/B 2.097720fF
C2 nand_0/A gnd! 6.253860fF
C3 nand_1/B gnd! 3.001320fF
C4 nand_1/A gnd! 6.522480fF
C5 nand_0/vdd gnd! 10.667521fF
C6 nand_0/gnd gnd! 8.607600fF
C7 S' gnd! 2.382240fF
C8 nand_2/vdd gnd! 8.912881fF
