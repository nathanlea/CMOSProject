magic
tech scmos
timestamp 1014240229
<< nwell >>
rect -4 26 25 83
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
<< ptransistor >>
rect 7 32 9 72
rect 12 32 14 72
<< ndiffusion >>
rect 6 6 7 16
rect 9 6 10 16
rect 14 6 15 16
rect 17 6 18 16
<< pdiffusion >>
rect 6 32 7 72
rect 9 32 12 72
rect 14 32 15 72
<< ndcontact >>
rect 2 6 6 16
rect 10 6 14 16
rect 18 6 22 16
<< pdcontact >>
rect 2 32 6 72
rect 15 32 19 72
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect 1 76 5 80
rect 14 76 18 80
<< polysilicon >>
rect 7 72 9 74
rect 12 72 14 74
rect 7 23 9 32
rect 6 19 9 23
rect 7 16 9 19
rect 12 29 14 32
rect 12 25 13 29
rect 12 19 14 25
rect 12 17 17 19
rect 15 16 17 17
rect 7 4 9 6
rect 15 4 17 6
<< polycontact >>
rect 2 19 6 23
rect 13 25 17 29
<< metal1 >>
rect -4 80 25 81
rect -4 76 1 80
rect 5 76 14 80
rect 18 76 25 80
rect -4 75 25 76
rect 2 72 6 75
rect 19 32 23 35
rect -4 26 13 29
rect -4 19 2 22
rect 20 22 23 32
rect 11 19 23 22
rect 11 16 14 19
rect 2 3 6 6
rect 18 3 22 6
rect -4 2 25 3
rect -4 -2 -2 2
rect 2 -2 14 2
rect 18 -2 25 2
rect -4 -3 25 -2
<< labels >>
rlabel metal1 9 0 9 0 8 gnd
rlabel metal1 -3 21 -3 21 3 A
rlabel metal1 22 28 22 28 7 Y
rlabel metal1 -3 27 -3 27 3 B
rlabel metal1 6 78 6 78 5 vdd
<< end >>
