* FILE: 21mux.sp

********************** begin header *****************************

* Sample Spice Header file for Generic 2.5V 0.25 um process (mmi25)

.OPTIONS post NOMOD post_version=9601

**################################################
* Only Typical/Typical spice models included
.include '${MMI_TOOLS}/sue/schematics/mspice/mmi25.mod'
* NOTE: these are contrived spice models
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=0,2,10,12 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3,13 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.6u
.param lp_min   =  0.6u

* used in source/drain area/perimeter calculation
.param sdd        =  0.66

.PARAM vddp=2.25	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "21mux" generated by MMI_SUE5.6.18 on Sun Nov 08 
*+ 19:54:31 CST 2015.

.SUBCKT nand2 in0 in1 out WP=2 WN=2
M_1 out in0 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_2 out in0 net_1 gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_3 out in1 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_4 net_1 in1 gnd gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
.ENDS	$ nand2

.SUBCKT inverter in out WP=2 LP=lp_min WN=1 LN=ln_min
M_1 out in gnd gnd n W='WN*1u' L=LN ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_2 out in vdd vdd p W='WP*1u' L=LP ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
.ENDS	$ inverter

* start main CELL 21mux
* .SUBCKT 21mux A B Out S 
Xnand2 B S net_3 nand2 
Xnand2_1 net_2 A net_1 nand2 
Xnand2_2 net_3 net_1 Out nand2 
Xinverter S net_2 inverter 
* .ENDS	$ 21mux

.GLOBAL gnd vdd

.END

