magic
tech scmos
timestamp 1447696045
<< nwell >>
rect -98 64 -13 75
rect -98 14 34 64
<< metal1 >>
rect -30 184 34 190
rect -56 145 -23 148
rect -56 138 -26 142
rect -96 120 -32 126
rect -36 112 -32 120
rect -36 100 34 112
rect -36 98 -24 100
rect -104 86 -88 89
rect -44 86 -36 90
rect -104 -28 -100 86
rect 32 71 42 74
rect -96 12 34 26
rect -104 -32 -68 -28
rect -103 -42 -77 -38
rect 8 -42 36 -38
rect -89 -52 -83 -48
rect 32 -73 36 -42
rect 32 -78 36 -77
rect -94 -97 32 -82
rect 39 -145 42 71
rect 10 -149 42 -145
rect -82 -198 18 -192
<< m2contact >>
rect 29 132 33 136
rect -36 86 -32 90
rect -92 76 -88 80
rect -107 -42 -103 -38
rect -93 -52 -89 -48
rect 32 -77 36 -73
<< metal2 >>
rect 33 132 43 136
rect -56 128 -32 131
rect -36 90 -32 128
rect -107 76 -92 80
rect -107 -38 -103 76
rect 39 23 43 132
rect -93 19 43 23
rect -93 -48 -89 19
rect 25 -61 47 -58
rect 32 -85 36 -77
rect -86 -89 36 -85
rect -86 -140 -82 -89
rect -30 -203 -26 -197
use ../../XOR2/magic/xor2  xor2_0 ../../XOR2/magic
timestamp 1160719867
transform -1 0 -23 0 -1 123
box 10 -3 75 105
use ../../mux21/magic/mux21  mux21_0 ../../mux21/magic
timestamp 1447275876
transform 1 0 -29 0 1 108
box -1 -90 63 84
use ../../FA/magic/fa  fa_0 ../../FA/magic
timestamp 1014102789
transform 1 0 -90 0 1 -85
box -5 -3 124 105
use ../../dffpos/magic/dffpos  dffpos_0 ../../dffpos/magic
timestamp 1447691457
transform 1 0 -44 0 -1 -184
box -38 -93 62 16
<< labels >>
rlabel metal1 1 186 1 186 1 vdd
rlabel metal1 -18 105 -18 105 1 gnd
rlabel metal1 -37 18 -37 18 1 vdd
rlabel metal1 -53 -90 -53 -90 1 gnd
rlabel metal2 -28 -202 -28 -202 1 clk
rlabel metal1 -24 -196 -24 -196 1 vdd
rlabel metal2 45 -60 45 -60 7 Cout
rlabel metal2 -54 129 -54 129 1 A
rlabel metal1 -55 146 -55 146 1 B
rlabel metal1 -102 88 -102 88 3 subtract
rlabel metal1 34 -40 34 -40 1 sum
rlabel metal1 -55 139 -55 139 1 S
rlabel metal2 -98 78 -98 78 1 Y
<< end >>
