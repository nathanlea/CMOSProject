magic
tech scmos
timestamp 1447439268
<< ntransistor >>
rect -29 -84 -27 -64
rect -21 -84 -19 -74
rect -16 -84 -14 -74
rect -7 -84 -5 -74
rect -2 -84 0 -74
rect 7 -84 9 -74
rect 23 -84 25 -74
rect 28 -84 30 -74
rect 38 -84 40 -74
rect 43 -84 45 -74
rect 51 -84 53 -64
<< ptransistor >>
rect -29 -35 -27 5
rect -21 -15 -19 5
rect -15 -15 -13 5
rect -7 -15 -5 5
rect -1 -15 1 5
rect 7 -15 9 5
rect 23 -15 25 5
rect 28 -15 30 5
rect 38 -5 40 5
rect 43 -5 45 5
rect 51 -35 53 5
<< ndiffusion >>
rect -30 -84 -29 -64
rect -27 -84 -26 -64
rect 46 -65 51 -64
rect -22 -84 -21 -74
rect -19 -84 -16 -74
rect -14 -84 -13 -74
rect -8 -84 -7 -74
rect -5 -84 -2 -74
rect 0 -84 1 -74
rect 6 -84 7 -74
rect 9 -84 10 -74
rect 22 -84 23 -74
rect 25 -84 28 -74
rect 30 -84 31 -74
rect 37 -84 38 -74
rect 40 -84 43 -74
rect 45 -84 46 -74
rect 50 -84 51 -65
rect 53 -84 54 -64
<< pdiffusion >>
rect -30 -35 -29 5
rect -27 -34 -26 5
rect -22 -15 -21 5
rect -19 -15 -15 5
rect -13 -15 -12 5
rect -8 -15 -7 5
rect -5 -15 -1 5
rect 1 -15 2 5
rect 6 -15 7 5
rect 9 -15 10 5
rect 22 -15 23 5
rect 25 -15 28 5
rect 30 -15 31 5
rect 37 -5 38 5
rect 40 -5 43 5
rect 45 -5 46 5
rect -27 -35 -22 -34
rect 50 -35 51 5
rect 53 -35 54 5
<< ndcontact >>
rect -34 -84 -30 -64
rect -26 -84 -22 -64
rect -13 -84 -8 -74
rect 1 -84 6 -74
rect 10 -84 14 -74
rect 18 -84 22 -74
rect 31 -84 37 -74
rect 46 -84 50 -65
rect 54 -84 58 -64
<< pdcontact >>
rect -34 -35 -30 5
rect -26 -34 -22 5
rect -12 -15 -8 5
rect 2 -15 6 5
rect 10 -15 14 5
rect 18 -15 22 5
rect 31 -15 37 5
rect 46 -35 50 5
rect 54 -35 58 5
<< psubstratepcontact >>
rect -38 -92 -34 -88
rect -21 -92 -17 -88
rect -6 -92 -2 -88
rect 10 -92 14 -88
rect 24 -92 28 -88
rect 42 -92 46 -88
<< nsubstratencontact >>
rect -38 9 -34 13
rect -21 9 -17 13
rect -5 9 -1 13
rect 10 9 14 13
rect 24 9 28 13
rect 43 9 47 13
<< polysilicon >>
rect -29 5 -27 7
rect -21 5 -19 7
rect -15 5 -13 7
rect -7 5 -5 7
rect -1 5 1 7
rect 7 5 9 7
rect 23 5 25 7
rect 28 5 30 7
rect 38 5 40 7
rect 43 5 45 7
rect 51 5 53 7
rect -29 -64 -27 -35
rect -21 -44 -19 -15
rect -21 -74 -19 -48
rect -15 -52 -13 -15
rect -7 -36 -5 -15
rect -7 -61 -5 -40
rect -16 -63 -5 -61
rect -1 -19 1 -15
rect -16 -74 -14 -63
rect -1 -66 1 -23
rect 7 -28 9 -15
rect 23 -17 25 -15
rect 14 -19 25 -17
rect -6 -71 -5 -67
rect -7 -74 -5 -71
rect -2 -70 -1 -66
rect -2 -74 0 -70
rect 7 -74 9 -32
rect 13 -71 15 -23
rect 28 -27 30 -15
rect 38 -22 40 -5
rect 36 -24 40 -22
rect 23 -29 30 -27
rect 21 -66 23 -57
rect 28 -59 30 -29
rect 43 -37 45 -5
rect 39 -39 45 -37
rect 38 -59 40 -43
rect 51 -45 53 -35
rect 49 -49 53 -45
rect 28 -61 35 -59
rect 21 -68 30 -66
rect 13 -73 25 -71
rect 23 -74 25 -73
rect 28 -74 30 -68
rect 33 -71 35 -61
rect 38 -63 39 -59
rect 33 -73 40 -71
rect 38 -74 40 -73
rect 43 -74 45 -59
rect 51 -64 53 -49
rect -29 -86 -27 -84
rect -21 -86 -19 -84
rect -16 -86 -14 -84
rect -7 -86 -5 -84
rect -2 -86 0 -84
rect 7 -86 9 -84
rect 23 -86 25 -84
rect 28 -86 30 -84
rect 38 -86 40 -84
rect 43 -86 45 -84
rect 51 -86 53 -84
<< polycontact >>
rect -33 -56 -29 -52
rect -23 -48 -19 -44
rect -9 -40 -5 -36
rect -15 -56 -11 -52
rect -1 -23 3 -19
rect 5 -32 9 -28
rect -10 -71 -6 -67
rect -1 -70 3 -66
rect 13 -23 17 -19
rect 19 -31 23 -27
rect 34 -28 38 -24
rect 19 -57 23 -53
rect 37 -43 41 -39
rect 45 -49 49 -45
rect 39 -63 43 -59
<< metal1 >>
rect -38 13 62 14
rect -34 9 -21 13
rect -17 9 -5 13
rect -1 9 10 13
rect 14 9 24 13
rect 28 9 43 13
rect 47 9 62 13
rect -38 8 62 9
rect -26 5 -22 8
rect 2 5 6 8
rect 18 5 22 8
rect 46 5 50 8
rect -18 -15 -12 -11
rect 30 -15 31 -10
rect 10 -19 13 -15
rect 3 -22 13 -19
rect -14 -32 5 -29
rect 12 -30 19 -27
rect 12 -36 15 -30
rect 31 -34 34 -24
rect -30 -39 -9 -37
rect -34 -40 -9 -39
rect -5 -39 15 -36
rect 22 -37 34 -34
rect -34 -41 -6 -40
rect -38 -47 -23 -44
rect -19 -47 2 -44
rect -29 -56 -15 -53
rect -11 -56 11 -53
rect 22 -53 25 -37
rect 41 -42 58 -39
rect 34 -49 45 -46
rect 15 -56 19 -53
rect -9 -67 -6 -56
rect 23 -56 58 -53
rect 43 -60 58 -59
rect 43 -62 54 -60
rect 3 -70 13 -67
rect 10 -74 13 -70
rect -18 -78 -13 -74
rect 30 -78 31 -74
rect -26 -87 -22 -84
rect 1 -87 6 -84
rect 18 -87 22 -84
rect 46 -87 50 -84
rect -38 -88 62 -87
rect -34 -92 -21 -88
rect -17 -92 -6 -88
rect -2 -92 10 -88
rect 14 -92 24 -88
rect 28 -92 42 -88
rect 46 -92 62 -88
rect -38 -93 62 -92
<< m2contact >>
rect -18 -19 -14 -15
rect 30 -19 34 -15
rect -18 -32 -14 -28
rect -34 -39 -30 -35
rect 11 -56 15 -52
rect 54 -39 58 -35
rect 30 -50 34 -46
rect -34 -64 -30 -60
rect 54 -64 58 -60
rect -18 -74 -14 -70
rect 30 -74 34 -70
<< metal2 >>
rect -18 -28 -14 -19
rect -34 -60 -30 -39
rect -18 -70 -14 -32
rect 14 -52 18 16
rect 15 -56 18 -52
rect 14 -93 18 -56
rect 30 -46 34 -19
rect 30 -70 34 -50
rect 54 -60 58 -39
<< labels >>
rlabel metal1 6 10 6 10 1 vdd
rlabel metal1 6 -91 6 -91 1 gnd
rlabel metal1 -37 -45 -37 -45 3 D
rlabel metal2 56 -48 56 -48 1 Q
rlabel metal2 16 15 16 15 5 clk
<< end >>
