magic
tech scmos
timestamp 1449155358
<< metal1 >>
rect -132 491 1451 503
rect -132 -135 -120 491
rect -108 467 1427 479
rect -108 329 -96 467
rect -83 387 1403 393
rect 25 351 29 379
rect 37 366 40 380
rect 25 348 58 351
rect -86 341 59 345
rect 159 341 163 359
rect 205 351 209 376
rect 224 363 228 376
rect 205 348 229 351
rect 209 341 224 345
rect 329 336 333 358
rect 374 351 378 378
rect 392 365 396 378
rect 374 348 396 351
rect 379 342 395 345
rect 499 338 503 350
rect 529 351 533 377
rect 548 364 552 377
rect 529 348 571 351
rect 533 342 566 345
rect 684 339 688 360
rect 712 351 716 379
rect 728 366 732 379
rect 712 348 733 351
rect 716 342 732 345
rect 856 338 859 364
rect 884 351 889 377
rect 899 365 904 377
rect 884 348 908 351
rect 888 341 908 344
rect 1023 339 1027 364
rect 1058 351 1062 377
rect 1074 364 1078 377
rect 1058 348 1082 351
rect 1187 339 1191 365
rect 1201 344 1204 348
rect 1225 348 1240 351
rect 1201 341 1240 344
rect -108 323 75 329
rect -108 121 -96 323
rect 71 315 75 323
rect 169 323 189 329
rect 340 323 357 329
rect 511 323 528 329
rect 672 323 701 329
rect 846 323 864 329
rect 1013 323 1034 329
rect 1177 323 1200 329
rect 169 315 179 323
rect 340 315 346 323
rect 511 315 516 323
rect 672 315 679 323
rect 71 303 179 315
rect 313 303 346 315
rect 482 303 516 315
rect 583 303 679 315
rect 846 315 851 323
rect 1013 316 1019 323
rect -6 289 -1 292
rect 3 289 8 292
rect 163 289 181 292
rect 333 289 346 292
rect 503 289 521 292
rect 684 289 688 312
rect 822 303 851 315
rect 856 289 859 306
rect 991 303 1019 316
rect 1177 315 1182 323
rect 1023 289 1027 313
rect 1158 303 1182 315
rect 1415 315 1427 467
rect 1187 289 1191 312
rect 1321 303 1427 315
rect -73 215 1398 229
rect -3 171 17 175
rect 165 171 184 175
rect 337 171 352 175
rect 507 171 520 175
rect 678 171 692 175
rect 847 171 859 175
rect 1009 171 1026 175
rect 1171 171 1191 175
rect 1009 142 1013 171
rect 1171 142 1175 171
rect 1319 156 1323 161
rect 1338 142 1342 145
rect 1415 121 1427 303
rect -108 106 1427 121
rect -108 -67 -96 106
rect -83 5 1403 11
rect -32 -34 -24 -31
rect 39 -34 43 -2
rect 14 -38 43 -34
rect -32 -41 -24 -38
rect -8 -47 3 -44
rect 0 -51 3 -47
rect 154 -60 158 -2
rect 326 -52 330 -5
rect 494 -45 499 -3
rect 666 -38 670 -2
rect 835 -31 839 -3
rect 1004 -24 1008 -3
rect 1171 -12 1175 -3
rect -108 -73 24 -67
rect -108 -111 -96 -73
rect 1415 -110 1427 106
rect 1277 -111 1427 -110
rect -108 -123 1427 -111
rect 1439 -134 1451 491
rect 1277 -135 1451 -134
rect -132 -147 1451 -135
rect 1439 -149 1451 -147
<< m2contact >>
rect -120 387 -115 393
rect -88 387 -83 393
rect 1403 387 1410 395
rect 25 379 29 383
rect 37 380 41 384
rect 205 376 209 380
rect 37 362 41 366
rect 159 359 163 363
rect -91 341 -86 345
rect 224 376 228 380
rect 224 359 228 363
rect 374 378 378 382
rect 329 358 333 362
rect 205 341 209 345
rect 159 337 163 341
rect 392 378 396 382
rect 392 361 396 365
rect 529 377 533 381
rect 499 350 503 354
rect 374 341 379 345
rect 329 332 333 336
rect 548 377 552 381
rect 712 379 716 383
rect 548 360 552 364
rect 684 360 688 364
rect 529 341 533 345
rect 499 334 503 338
rect 728 379 732 383
rect 884 377 889 382
rect 728 362 732 366
rect 856 364 860 368
rect 712 341 716 345
rect 684 334 689 339
rect 899 377 904 382
rect 1058 377 1062 381
rect 899 360 904 365
rect 1023 364 1028 369
rect 884 341 888 345
rect 1074 377 1078 381
rect 1074 360 1078 364
rect 1187 365 1192 370
rect 1064 341 1068 345
rect 1201 348 1205 352
rect 1220 347 1225 351
rect 856 334 860 338
rect 1023 334 1028 339
rect 1187 334 1192 339
rect -120 215 -112 223
rect 684 312 689 317
rect -1 289 3 293
rect 159 289 163 293
rect 329 289 333 293
rect 499 289 503 293
rect 856 306 860 310
rect 1023 313 1028 318
rect 1187 312 1192 317
rect 1432 387 1439 395
rect -85 215 -73 229
rect 1398 215 1411 229
rect -9 171 -3 177
rect 161 171 165 175
rect 333 171 337 175
rect 503 171 507 175
rect 674 171 678 175
rect 842 171 847 176
rect 161 142 166 147
rect 333 142 338 147
rect 503 142 508 147
rect 674 142 679 147
rect 842 142 847 147
rect 1431 215 1439 223
rect -120 5 -112 14
rect -91 5 -83 14
rect 1403 5 1409 12
rect 39 -2 43 2
rect 154 -2 158 2
rect 326 -5 330 -1
rect 494 -3 499 2
rect 666 -2 670 2
rect 835 -3 839 1
rect 1004 -3 1008 1
rect 1171 -3 1175 1
rect 1171 -17 1176 -12
rect 1008 -24 1012 -20
rect 839 -31 844 -26
rect 670 -38 675 -33
rect 499 -45 504 -40
rect 330 -52 335 -47
rect 158 -60 164 -54
rect 1433 5 1439 12
<< metal2 >>
rect -115 387 -88 392
rect 25 383 28 511
rect 37 384 40 511
rect 205 397 208 511
rect 224 397 227 511
rect 205 380 209 397
rect 224 380 228 397
rect 374 396 377 511
rect 392 396 395 511
rect 529 396 532 511
rect 548 396 551 511
rect 374 382 378 396
rect 392 382 396 396
rect 529 381 533 396
rect 548 381 552 396
rect 712 395 715 511
rect 728 395 731 511
rect 884 396 887 511
rect 899 396 902 511
rect 1058 396 1061 511
rect 1074 396 1077 511
rect 1220 396 1223 511
rect 1231 396 1234 511
rect 712 383 716 395
rect 728 383 732 395
rect 884 382 889 396
rect 899 382 904 396
rect 1058 381 1062 396
rect 1074 381 1078 396
rect -1 370 1192 372
rect -1 369 1187 370
rect -139 341 -91 345
rect -1 293 3 369
rect 159 363 163 369
rect 37 334 40 362
rect 98 348 186 351
rect 98 341 101 348
rect 183 345 186 348
rect 183 341 205 345
rect 37 331 58 334
rect 159 293 163 337
rect 224 331 228 359
rect 329 362 333 369
rect 270 348 366 352
rect 270 341 274 348
rect 362 345 366 348
rect 362 341 374 345
rect 329 293 333 332
rect 392 331 396 361
rect 499 354 502 369
rect 684 364 688 369
rect 856 368 860 369
rect 439 349 478 352
rect 439 341 443 349
rect 475 345 478 349
rect 475 342 529 345
rect 548 334 552 360
rect 613 349 686 352
rect 613 341 616 349
rect 683 345 686 349
rect 683 342 712 345
rect 499 293 502 334
rect 548 331 571 334
rect 684 317 689 334
rect 728 334 732 362
rect 782 351 852 352
rect 782 348 866 351
rect 782 341 786 348
rect 863 344 866 348
rect 863 341 884 344
rect 899 334 904 360
rect 951 348 1043 352
rect 951 341 955 348
rect 1039 345 1043 348
rect 1039 341 1064 345
rect 1074 334 1078 360
rect 1118 348 1201 351
rect 1220 351 1225 396
rect 1118 341 1122 348
rect 1231 334 1236 396
rect 1410 387 1432 393
rect 728 331 734 334
rect 856 310 859 334
rect 899 331 908 334
rect 1023 318 1027 334
rect 1074 331 1082 334
rect 1187 317 1191 334
rect 1231 331 1239 334
rect -9 286 3 289
rect -112 215 -85 223
rect -9 177 -5 286
rect 1411 215 1431 223
rect 161 147 165 171
rect 333 147 337 171
rect 503 147 506 171
rect 674 147 678 171
rect 842 147 846 171
rect 150 142 151 145
rect 322 142 323 145
rect 662 142 663 145
rect -112 5 -91 11
rect 77 1 150 3
rect 43 0 150 1
rect 43 -2 81 0
rect 147 -7 150 0
rect 154 2 158 65
rect 161 0 322 3
rect 161 -7 164 0
rect 147 -10 164 -7
rect 319 -8 322 0
rect 326 -1 330 62
rect 334 0 491 3
rect 334 -8 337 0
rect 319 -11 337 -8
rect 488 -7 491 0
rect 494 2 499 63
rect 811 62 812 65
rect 967 62 970 65
rect 502 0 663 3
rect 502 -7 505 0
rect 488 -10 505 -7
rect 660 -5 663 0
rect 666 2 670 62
rect 673 0 831 3
rect 673 -5 676 0
rect 660 -8 676 -5
rect 827 -6 831 0
rect 835 1 839 62
rect 843 0 1000 3
rect 843 -6 846 0
rect 827 -9 846 -6
rect 996 -6 1000 0
rect 1004 1 1008 62
rect 1012 0 1167 3
rect 1012 -6 1016 0
rect 996 -9 1016 -6
rect 1163 -6 1167 0
rect 1171 1 1175 63
rect 1249 62 1254 65
rect 1334 3 1338 65
rect 1409 5 1433 11
rect 1179 0 1261 3
rect 1179 -6 1182 0
rect 1163 -9 1182 -6
rect 1333 -6 1338 3
rect 1333 -10 1492 -6
rect 1176 -17 1492 -13
rect 1012 -24 1492 -20
rect 844 -31 1492 -27
rect 675 -38 1492 -34
rect 504 -45 1492 -41
rect 335 -52 1492 -48
rect 164 -60 1492 -55
use ../../nand/magic/nand  nand_0 ../../nand/magic
timestamp 1013989602
transform 1 0 -28 0 1 -70
box -4 -3 28 83
use ../../bitslice/magic/bitslice  bitslice_0 ../../bitslice/magic
timestamp 1449109615
transform 1 0 107 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_1
timestamp 1449109615
transform 1 0 279 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_2
timestamp 1449109615
transform 1 0 448 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_3
timestamp 1449109615
transform 1 0 619 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_4
timestamp 1449109615
transform 1 0 788 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_5
timestamp 1449109615
transform 1 0 957 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_6
timestamp 1449109615
transform 1 0 1124 0 1 203
box -107 -203 55 192
use ../../bitslice/magic/bitslice  bitslice_7
timestamp 1449109615
transform 1 0 1287 0 1 203
box -107 -203 55 192
use ../../inv/magic/inverter  inverter_0 ../../inv/magic
timestamp 1013989724
transform 1 0 4 0 1 -72
box -4 -1 20 85
<< labels >>
rlabel metal1 -28 -33 -28 -33 3 clk
rlabel metal1 -29 -40 -29 -40 3 loadR
rlabel metal1 -4 291 -4 291 1 subtract
rlabel metal2 1251 64 1251 64 1 Out7
rlabel metal1 1341 144 1341 144 7 Cout
rlabel metal1 1321 158 1321 158 1 gundy
rlabel metal1 -126 497 -126 497 1 Vdd
rlabel metal1 -101 471 -101 471 1 Gnd
rlabel metal2 1490 -8 1490 -8 7 Out7
rlabel metal2 1490 -15 1490 -15 7 Out6
rlabel metal2 1490 -22 1490 -22 7 Out5
rlabel metal2 1490 -29 1490 -29 7 Out4
rlabel metal2 1490 -36 1490 -36 7 Out3
rlabel metal2 1490 -43 1490 -43 7 Out2
rlabel metal2 1490 -50 1490 -50 7 Out1
rlabel metal2 1490 -58 1490 -58 7 Out0
rlabel metal2 -137 343 -137 343 3 loadB
rlabel metal2 26 509 26 509 5 B0
rlabel metal2 38 509 38 509 5 A0
rlabel metal2 206 509 206 509 5 B1
rlabel metal2 225 509 225 509 5 A1
rlabel metal2 375 509 375 509 5 B2
rlabel metal2 393 509 393 509 5 A2
rlabel metal2 530 509 530 509 5 B3
rlabel metal2 549 509 549 509 5 A3
rlabel metal2 713 509 713 509 5 B4
rlabel metal2 729 509 729 509 5 A4
rlabel metal2 885 508 885 508 5 B5
rlabel metal2 900 508 900 508 5 A5
rlabel metal2 1059 508 1059 508 5 B6
rlabel metal2 1075 508 1075 508 5 A6
rlabel metal2 1221 508 1221 508 5 B7
rlabel metal2 1232 508 1232 508 5 A7
<< end >>
