* SPICE3 file created from prjMagic.ext - technology: scmos

.option scale=0.3u

M1000 inverter_0/Y inverter_0/A Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=20220 ps=8806
M1001 inverter_0/Y inverter_0/A Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=10230 ps=4992
M1002 Vdd inverter_0/Y bitslice_7/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1003 bitslice_7/dffpos_0/a_n19_n15# gundy Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1004 bitslice_7/dffpos_0/a_n14_n84# inverter_0/Y bitslice_7/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1005 bitslice_7/dffpos_0/a_n5_n15# bitslice_7/dffpos_0/a_n34_n84# bitslice_7/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1006 Vdd bitslice_7/dffpos_0/a_n2_n86# bitslice_7/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 bitslice_7/dffpos_0/a_n2_n86# bitslice_7/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1008 bitslice_7/dffpos_0/a_25_n15# bitslice_7/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1009 bitslice_7/dffpos_0/a_30_n84# bitslice_7/dffpos_0/a_n34_n84# bitslice_7/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1010 bitslice_7/dffpos_0/a_40_n5# inverter_0/Y bitslice_7/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1011 Vdd Out7 bitslice_7/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 Gnd inverter_0/Y bitslice_7/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1013 Out7 bitslice_7/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1014 bitslice_7/dffpos_0/a_n19_n84# gundy Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1015 bitslice_7/dffpos_0/a_n14_n84# bitslice_7/dffpos_0/a_n34_n84# bitslice_7/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1016 bitslice_7/dffpos_0/a_n5_n84# inverter_0/Y bitslice_7/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1017 Gnd bitslice_7/dffpos_0/a_n2_n86# bitslice_7/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1018 bitslice_7/dffpos_0/a_n2_n86# bitslice_7/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1019 bitslice_7/dffpos_0/a_25_n84# bitslice_7/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1020 bitslice_7/dffpos_0/a_30_n84# inverter_0/Y bitslice_7/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1021 bitslice_7/dffpos_0/a_40_n84# bitslice_7/dffpos_0/a_n34_n84# bitslice_7/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1022 Gnd Out7 bitslice_7/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 Out7 bitslice_7/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1024 Vdd bitslice_7/fa_0/A bitslice_7/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1025 bitslice_7/fa_0/a_2_74# bitslice_7/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 bitslice_7/fa_0/a_25_6# bitslice_7/Cin bitslice_7/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1027 bitslice_7/fa_0/a_33_74# bitslice_7/Y bitslice_7/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1028 Vdd bitslice_7/fa_0/A bitslice_7/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1029 bitslice_7/fa_0/a_46_74# bitslice_7/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1030 Vdd bitslice_7/Y bitslice_7/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1031 bitslice_7/fa_0/a_46_74# bitslice_7/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 bitslice_7/fa_0/a_70_6# bitslice_7/fa_0/a_25_6# bitslice_7/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1033 bitslice_7/fa_0/a_79_74# bitslice_7/Cin bitslice_7/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1034 bitslice_7/fa_0/a_84_74# bitslice_7/Y bitslice_7/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1035 Vdd bitslice_7/fa_0/A bitslice_7/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 gundy bitslice_7/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1037 Cout bitslice_7/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1038 Gnd bitslice_7/fa_0/A bitslice_7/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1039 bitslice_7/fa_0/a_2_6# bitslice_7/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 bitslice_7/fa_0/a_25_6# bitslice_7/Cin bitslice_7/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1041 bitslice_7/fa_0/a_33_6# bitslice_7/Y bitslice_7/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1042 Gnd bitslice_7/fa_0/A bitslice_7/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 bitslice_7/fa_0/a_46_6# bitslice_7/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1044 Gnd bitslice_7/Y bitslice_7/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 bitslice_7/fa_0/a_46_6# bitslice_7/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1046 bitslice_7/fa_0/a_70_6# bitslice_7/fa_0/a_25_6# bitslice_7/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1047 bitslice_7/fa_0/a_79_6# bitslice_7/Cin bitslice_7/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1048 bitslice_7/fa_0/a_84_6# bitslice_7/Y bitslice_7/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1049 Gnd bitslice_7/fa_0/A bitslice_7/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 gundy bitslice_7/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1051 Cout bitslice_7/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1052 bitslice_7/mux21_0/nand_1/A Out7 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1053 Vdd bitslice_7/mux21_0/nand_2/B bitslice_7/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 bitslice_7/mux21_0/nand_2/a_9_6# Out7 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1055 bitslice_7/mux21_0/nand_1/A bitslice_7/mux21_0/nand_2/B bitslice_7/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1056 bitslice_7/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1057 bitslice_7/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1058 bitslice_7/fa_0/A bitslice_7/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1059 Vdd bitslice_7/mux21_0/nand_1/B bitslice_7/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 bitslice_7/mux21_0/nand_1/a_9_6# bitslice_7/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1061 bitslice_7/fa_0/A bitslice_7/mux21_0/nand_1/B bitslice_7/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1062 bitslice_7/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1063 Vdd B7 bitslice_7/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 bitslice_7/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1065 bitslice_7/mux21_0/nand_1/B B7 bitslice_7/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1066 Vdd A7 bitslice_7/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1067 bitslice_7/xor2_0/a_33_54# bitslice_7/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1068 bitslice_7/Y A7 bitslice_7/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1069 bitslice_7/xor2_0/a_50_54# bitslice_7/xor2_0/a_17_6# bitslice_7/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1070 Vdd subtract bitslice_7/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1071 bitslice_7/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1072 Gnd A7 bitslice_7/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1073 bitslice_7/xor2_0/a_33_6# bitslice_7/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1074 bitslice_7/Y bitslice_7/xor2_0/a_17_6# bitslice_7/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1075 bitslice_7/xor2_0/a_50_6# A7 bitslice_7/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1076 Gnd subtract bitslice_7/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1077 bitslice_7/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1078 Vdd inverter_0/Y bitslice_6/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1079 bitslice_6/dffpos_0/a_n19_n15# bitslice_6/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1080 bitslice_6/dffpos_0/a_n14_n84# inverter_0/Y bitslice_6/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1081 bitslice_6/dffpos_0/a_n5_n15# bitslice_6/dffpos_0/a_n34_n84# bitslice_6/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1082 Vdd bitslice_6/dffpos_0/a_n2_n86# bitslice_6/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 bitslice_6/dffpos_0/a_n2_n86# bitslice_6/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1084 bitslice_6/dffpos_0/a_25_n15# bitslice_6/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1085 bitslice_6/dffpos_0/a_30_n84# bitslice_6/dffpos_0/a_n34_n84# bitslice_6/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1086 bitslice_6/dffpos_0/a_40_n5# inverter_0/Y bitslice_6/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1087 Vdd Out6 bitslice_6/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 Gnd inverter_0/Y bitslice_6/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1089 Out6 bitslice_6/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1090 bitslice_6/dffpos_0/a_n19_n84# bitslice_6/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1091 bitslice_6/dffpos_0/a_n14_n84# bitslice_6/dffpos_0/a_n34_n84# bitslice_6/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1092 bitslice_6/dffpos_0/a_n5_n84# inverter_0/Y bitslice_6/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1093 Gnd bitslice_6/dffpos_0/a_n2_n86# bitslice_6/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 bitslice_6/dffpos_0/a_n2_n86# bitslice_6/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1095 bitslice_6/dffpos_0/a_25_n84# bitslice_6/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1096 bitslice_6/dffpos_0/a_30_n84# inverter_0/Y bitslice_6/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1097 bitslice_6/dffpos_0/a_40_n84# bitslice_6/dffpos_0/a_n34_n84# bitslice_6/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1098 Gnd Out6 bitslice_6/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1099 Out6 bitslice_6/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1100 Vdd bitslice_6/fa_0/A bitslice_6/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1101 bitslice_6/fa_0/a_2_74# bitslice_6/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 bitslice_6/fa_0/a_25_6# bitslice_6/Cin bitslice_6/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1103 bitslice_6/fa_0/a_33_74# bitslice_6/Y bitslice_6/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1104 Vdd bitslice_6/fa_0/A bitslice_6/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1105 bitslice_6/fa_0/a_46_74# bitslice_6/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1106 Vdd bitslice_6/Y bitslice_6/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 bitslice_6/fa_0/a_46_74# bitslice_6/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 bitslice_6/fa_0/a_70_6# bitslice_6/fa_0/a_25_6# bitslice_6/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1109 bitslice_6/fa_0/a_79_74# bitslice_6/Cin bitslice_6/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1110 bitslice_6/fa_0/a_84_74# bitslice_6/Y bitslice_6/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1111 Vdd bitslice_6/fa_0/A bitslice_6/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 bitslice_6/sum bitslice_6/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1113 bitslice_7/Cin bitslice_6/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1114 Gnd bitslice_6/fa_0/A bitslice_6/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1115 bitslice_6/fa_0/a_2_6# bitslice_6/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 bitslice_6/fa_0/a_25_6# bitslice_6/Cin bitslice_6/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1117 bitslice_6/fa_0/a_33_6# bitslice_6/Y bitslice_6/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1118 Gnd bitslice_6/fa_0/A bitslice_6/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 bitslice_6/fa_0/a_46_6# bitslice_6/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1120 Gnd bitslice_6/Y bitslice_6/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 bitslice_6/fa_0/a_46_6# bitslice_6/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 bitslice_6/fa_0/a_70_6# bitslice_6/fa_0/a_25_6# bitslice_6/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1123 bitslice_6/fa_0/a_79_6# bitslice_6/Cin bitslice_6/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1124 bitslice_6/fa_0/a_84_6# bitslice_6/Y bitslice_6/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1125 Gnd bitslice_6/fa_0/A bitslice_6/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 bitslice_6/sum bitslice_6/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1127 bitslice_7/Cin bitslice_6/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1128 bitslice_6/mux21_0/nand_1/A Out6 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1129 Vdd bitslice_6/mux21_0/nand_2/B bitslice_6/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 bitslice_6/mux21_0/nand_2/a_9_6# Out6 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1131 bitslice_6/mux21_0/nand_1/A bitslice_6/mux21_0/nand_2/B bitslice_6/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1132 bitslice_6/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1133 bitslice_6/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1134 bitslice_6/fa_0/A bitslice_6/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1135 Vdd bitslice_6/mux21_0/nand_1/B bitslice_6/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 bitslice_6/mux21_0/nand_1/a_9_6# bitslice_6/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1137 bitslice_6/fa_0/A bitslice_6/mux21_0/nand_1/B bitslice_6/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1138 bitslice_6/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1139 Vdd B6 bitslice_6/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 bitslice_6/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1141 bitslice_6/mux21_0/nand_1/B B6 bitslice_6/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1142 Vdd A6 bitslice_6/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1143 bitslice_6/xor2_0/a_33_54# bitslice_6/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1144 bitslice_6/Y A6 bitslice_6/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1145 bitslice_6/xor2_0/a_50_54# bitslice_6/xor2_0/a_17_6# bitslice_6/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1146 Vdd subtract bitslice_6/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 bitslice_6/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1148 Gnd A6 bitslice_6/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1149 bitslice_6/xor2_0/a_33_6# bitslice_6/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1150 bitslice_6/Y bitslice_6/xor2_0/a_17_6# bitslice_6/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1151 bitslice_6/xor2_0/a_50_6# A6 bitslice_6/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1152 Gnd subtract bitslice_6/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 bitslice_6/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1154 Vdd inverter_0/Y bitslice_5/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1155 bitslice_5/dffpos_0/a_n19_n15# bitslice_5/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1156 bitslice_5/dffpos_0/a_n14_n84# inverter_0/Y bitslice_5/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1157 bitslice_5/dffpos_0/a_n5_n15# bitslice_5/dffpos_0/a_n34_n84# bitslice_5/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1158 Vdd bitslice_5/dffpos_0/a_n2_n86# bitslice_5/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 bitslice_5/dffpos_0/a_n2_n86# bitslice_5/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1160 bitslice_5/dffpos_0/a_25_n15# bitslice_5/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1161 bitslice_5/dffpos_0/a_30_n84# bitslice_5/dffpos_0/a_n34_n84# bitslice_5/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1162 bitslice_5/dffpos_0/a_40_n5# inverter_0/Y bitslice_5/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1163 Vdd Out5 bitslice_5/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 Gnd inverter_0/Y bitslice_5/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1165 Out5 bitslice_5/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1166 bitslice_5/dffpos_0/a_n19_n84# bitslice_5/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1167 bitslice_5/dffpos_0/a_n14_n84# bitslice_5/dffpos_0/a_n34_n84# bitslice_5/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1168 bitslice_5/dffpos_0/a_n5_n84# inverter_0/Y bitslice_5/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1169 Gnd bitslice_5/dffpos_0/a_n2_n86# bitslice_5/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 bitslice_5/dffpos_0/a_n2_n86# bitslice_5/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1171 bitslice_5/dffpos_0/a_25_n84# bitslice_5/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1172 bitslice_5/dffpos_0/a_30_n84# inverter_0/Y bitslice_5/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1173 bitslice_5/dffpos_0/a_40_n84# bitslice_5/dffpos_0/a_n34_n84# bitslice_5/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1174 Gnd Out5 bitslice_5/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 Out5 bitslice_5/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1176 Vdd bitslice_5/fa_0/A bitslice_5/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1177 bitslice_5/fa_0/a_2_74# bitslice_5/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 bitslice_5/fa_0/a_25_6# bitslice_5/Cin bitslice_5/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1179 bitslice_5/fa_0/a_33_74# bitslice_5/Y bitslice_5/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1180 Vdd bitslice_5/fa_0/A bitslice_5/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 bitslice_5/fa_0/a_46_74# bitslice_5/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1182 Vdd bitslice_5/Y bitslice_5/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 bitslice_5/fa_0/a_46_74# bitslice_5/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 bitslice_5/fa_0/a_70_6# bitslice_5/fa_0/a_25_6# bitslice_5/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1185 bitslice_5/fa_0/a_79_74# bitslice_5/Cin bitslice_5/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1186 bitslice_5/fa_0/a_84_74# bitslice_5/Y bitslice_5/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1187 Vdd bitslice_5/fa_0/A bitslice_5/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 bitslice_5/sum bitslice_5/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1189 bitslice_6/Cin bitslice_5/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1190 Gnd bitslice_5/fa_0/A bitslice_5/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1191 bitslice_5/fa_0/a_2_6# bitslice_5/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 bitslice_5/fa_0/a_25_6# bitslice_5/Cin bitslice_5/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1193 bitslice_5/fa_0/a_33_6# bitslice_5/Y bitslice_5/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1194 Gnd bitslice_5/fa_0/A bitslice_5/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 bitslice_5/fa_0/a_46_6# bitslice_5/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1196 Gnd bitslice_5/Y bitslice_5/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 bitslice_5/fa_0/a_46_6# bitslice_5/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 bitslice_5/fa_0/a_70_6# bitslice_5/fa_0/a_25_6# bitslice_5/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1199 bitslice_5/fa_0/a_79_6# bitslice_5/Cin bitslice_5/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1200 bitslice_5/fa_0/a_84_6# bitslice_5/Y bitslice_5/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1201 Gnd bitslice_5/fa_0/A bitslice_5/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1202 bitslice_5/sum bitslice_5/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1203 bitslice_6/Cin bitslice_5/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1204 bitslice_5/mux21_0/nand_1/A Out5 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1205 Vdd bitslice_5/mux21_0/nand_2/B bitslice_5/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 bitslice_5/mux21_0/nand_2/a_9_6# Out5 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1207 bitslice_5/mux21_0/nand_1/A bitslice_5/mux21_0/nand_2/B bitslice_5/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1208 bitslice_5/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1209 bitslice_5/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1210 bitslice_5/fa_0/A bitslice_5/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1211 Vdd bitslice_5/mux21_0/nand_1/B bitslice_5/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 bitslice_5/mux21_0/nand_1/a_9_6# bitslice_5/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1213 bitslice_5/fa_0/A bitslice_5/mux21_0/nand_1/B bitslice_5/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1214 bitslice_5/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1215 Vdd B5 bitslice_5/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 bitslice_5/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1217 bitslice_5/mux21_0/nand_1/B B5 bitslice_5/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1218 Vdd A5 bitslice_5/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1219 bitslice_5/xor2_0/a_33_54# bitslice_5/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1220 bitslice_5/Y A5 bitslice_5/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1221 bitslice_5/xor2_0/a_50_54# bitslice_5/xor2_0/a_17_6# bitslice_5/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1222 Vdd subtract bitslice_5/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 bitslice_5/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1224 Gnd A5 bitslice_5/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1225 bitslice_5/xor2_0/a_33_6# bitslice_5/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1226 bitslice_5/Y bitslice_5/xor2_0/a_17_6# bitslice_5/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1227 bitslice_5/xor2_0/a_50_6# A5 bitslice_5/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1228 Gnd subtract bitslice_5/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 bitslice_5/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1230 Vdd inverter_0/Y bitslice_4/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1231 bitslice_4/dffpos_0/a_n19_n15# bitslice_4/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1232 bitslice_4/dffpos_0/a_n14_n84# inverter_0/Y bitslice_4/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1233 bitslice_4/dffpos_0/a_n5_n15# bitslice_4/dffpos_0/a_n34_n84# bitslice_4/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1234 Vdd bitslice_4/dffpos_0/a_n2_n86# bitslice_4/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 bitslice_4/dffpos_0/a_n2_n86# bitslice_4/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1236 bitslice_4/dffpos_0/a_25_n15# bitslice_4/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1237 bitslice_4/dffpos_0/a_30_n84# bitslice_4/dffpos_0/a_n34_n84# bitslice_4/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1238 bitslice_4/dffpos_0/a_40_n5# inverter_0/Y bitslice_4/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1239 Vdd Out4 bitslice_4/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 Gnd inverter_0/Y bitslice_4/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1241 Out4 bitslice_4/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1242 bitslice_4/dffpos_0/a_n19_n84# bitslice_4/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1243 bitslice_4/dffpos_0/a_n14_n84# bitslice_4/dffpos_0/a_n34_n84# bitslice_4/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1244 bitslice_4/dffpos_0/a_n5_n84# inverter_0/Y bitslice_4/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1245 Gnd bitslice_4/dffpos_0/a_n2_n86# bitslice_4/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 bitslice_4/dffpos_0/a_n2_n86# bitslice_4/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1247 bitslice_4/dffpos_0/a_25_n84# bitslice_4/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1248 bitslice_4/dffpos_0/a_30_n84# inverter_0/Y bitslice_4/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1249 bitslice_4/dffpos_0/a_40_n84# bitslice_4/dffpos_0/a_n34_n84# bitslice_4/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1250 Gnd Out4 bitslice_4/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 Out4 bitslice_4/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1252 Vdd bitslice_4/fa_0/A bitslice_4/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1253 bitslice_4/fa_0/a_2_74# bitslice_4/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1254 bitslice_4/fa_0/a_25_6# bitslice_4/Cin bitslice_4/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1255 bitslice_4/fa_0/a_33_74# bitslice_4/Y bitslice_4/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1256 Vdd bitslice_4/fa_0/A bitslice_4/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 bitslice_4/fa_0/a_46_74# bitslice_4/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1258 Vdd bitslice_4/Y bitslice_4/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 bitslice_4/fa_0/a_46_74# bitslice_4/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 bitslice_4/fa_0/a_70_6# bitslice_4/fa_0/a_25_6# bitslice_4/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1261 bitslice_4/fa_0/a_79_74# bitslice_4/Cin bitslice_4/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1262 bitslice_4/fa_0/a_84_74# bitslice_4/Y bitslice_4/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1263 Vdd bitslice_4/fa_0/A bitslice_4/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1264 bitslice_4/sum bitslice_4/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1265 bitslice_5/Cin bitslice_4/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1266 Gnd bitslice_4/fa_0/A bitslice_4/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1267 bitslice_4/fa_0/a_2_6# bitslice_4/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 bitslice_4/fa_0/a_25_6# bitslice_4/Cin bitslice_4/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1269 bitslice_4/fa_0/a_33_6# bitslice_4/Y bitslice_4/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1270 Gnd bitslice_4/fa_0/A bitslice_4/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 bitslice_4/fa_0/a_46_6# bitslice_4/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1272 Gnd bitslice_4/Y bitslice_4/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 bitslice_4/fa_0/a_46_6# bitslice_4/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 bitslice_4/fa_0/a_70_6# bitslice_4/fa_0/a_25_6# bitslice_4/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1275 bitslice_4/fa_0/a_79_6# bitslice_4/Cin bitslice_4/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1276 bitslice_4/fa_0/a_84_6# bitslice_4/Y bitslice_4/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1277 Gnd bitslice_4/fa_0/A bitslice_4/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1278 bitslice_4/sum bitslice_4/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1279 bitslice_5/Cin bitslice_4/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1280 bitslice_4/mux21_0/nand_1/A Out4 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1281 Vdd bitslice_4/mux21_0/nand_2/B bitslice_4/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 bitslice_4/mux21_0/nand_2/a_9_6# Out4 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1283 bitslice_4/mux21_0/nand_1/A bitslice_4/mux21_0/nand_2/B bitslice_4/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1284 bitslice_4/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1285 bitslice_4/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1286 bitslice_4/fa_0/A bitslice_4/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1287 Vdd bitslice_4/mux21_0/nand_1/B bitslice_4/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1288 bitslice_4/mux21_0/nand_1/a_9_6# bitslice_4/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1289 bitslice_4/fa_0/A bitslice_4/mux21_0/nand_1/B bitslice_4/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1290 bitslice_4/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1291 Vdd B4 bitslice_4/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 bitslice_4/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1293 bitslice_4/mux21_0/nand_1/B B4 bitslice_4/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1294 Vdd A4 bitslice_4/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1295 bitslice_4/xor2_0/a_33_54# bitslice_4/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1296 bitslice_4/Y A4 bitslice_4/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1297 bitslice_4/xor2_0/a_50_54# bitslice_4/xor2_0/a_17_6# bitslice_4/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1298 Vdd subtract bitslice_4/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 bitslice_4/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1300 Gnd A4 bitslice_4/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1301 bitslice_4/xor2_0/a_33_6# bitslice_4/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1302 bitslice_4/Y bitslice_4/xor2_0/a_17_6# bitslice_4/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1303 bitslice_4/xor2_0/a_50_6# A4 bitslice_4/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1304 Gnd subtract bitslice_4/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1305 bitslice_4/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1306 Vdd inverter_0/Y bitslice_3/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1307 bitslice_3/dffpos_0/a_n19_n15# bitslice_3/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1308 bitslice_3/dffpos_0/a_n14_n84# inverter_0/Y bitslice_3/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1309 bitslice_3/dffpos_0/a_n5_n15# bitslice_3/dffpos_0/a_n34_n84# bitslice_3/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1310 Vdd bitslice_3/dffpos_0/a_n2_n86# bitslice_3/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 bitslice_3/dffpos_0/a_n2_n86# bitslice_3/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1312 bitslice_3/dffpos_0/a_25_n15# bitslice_3/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1313 bitslice_3/dffpos_0/a_30_n84# bitslice_3/dffpos_0/a_n34_n84# bitslice_3/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1314 bitslice_3/dffpos_0/a_40_n5# inverter_0/Y bitslice_3/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1315 Vdd Out3 bitslice_3/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 Gnd inverter_0/Y bitslice_3/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1317 Out3 bitslice_3/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1318 bitslice_3/dffpos_0/a_n19_n84# bitslice_3/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1319 bitslice_3/dffpos_0/a_n14_n84# bitslice_3/dffpos_0/a_n34_n84# bitslice_3/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1320 bitslice_3/dffpos_0/a_n5_n84# inverter_0/Y bitslice_3/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1321 Gnd bitslice_3/dffpos_0/a_n2_n86# bitslice_3/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 bitslice_3/dffpos_0/a_n2_n86# bitslice_3/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1323 bitslice_3/dffpos_0/a_25_n84# bitslice_3/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1324 bitslice_3/dffpos_0/a_30_n84# inverter_0/Y bitslice_3/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1325 bitslice_3/dffpos_0/a_40_n84# bitslice_3/dffpos_0/a_n34_n84# bitslice_3/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1326 Gnd Out3 bitslice_3/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1327 Out3 bitslice_3/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1328 Vdd bitslice_3/fa_0/A bitslice_3/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1329 bitslice_3/fa_0/a_2_74# bitslice_3/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 bitslice_3/fa_0/a_25_6# bitslice_3/Cin bitslice_3/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1331 bitslice_3/fa_0/a_33_74# bitslice_3/Y bitslice_3/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1332 Vdd bitslice_3/fa_0/A bitslice_3/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 bitslice_3/fa_0/a_46_74# bitslice_3/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1334 Vdd bitslice_3/Y bitslice_3/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 bitslice_3/fa_0/a_46_74# bitslice_3/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 bitslice_3/fa_0/a_70_6# bitslice_3/fa_0/a_25_6# bitslice_3/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1337 bitslice_3/fa_0/a_79_74# bitslice_3/Cin bitslice_3/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1338 bitslice_3/fa_0/a_84_74# bitslice_3/Y bitslice_3/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1339 Vdd bitslice_3/fa_0/A bitslice_3/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 bitslice_3/sum bitslice_3/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1341 bitslice_4/Cin bitslice_3/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1342 Gnd bitslice_3/fa_0/A bitslice_3/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1343 bitslice_3/fa_0/a_2_6# bitslice_3/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1344 bitslice_3/fa_0/a_25_6# bitslice_3/Cin bitslice_3/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1345 bitslice_3/fa_0/a_33_6# bitslice_3/Y bitslice_3/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1346 Gnd bitslice_3/fa_0/A bitslice_3/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1347 bitslice_3/fa_0/a_46_6# bitslice_3/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1348 Gnd bitslice_3/Y bitslice_3/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1349 bitslice_3/fa_0/a_46_6# bitslice_3/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1350 bitslice_3/fa_0/a_70_6# bitslice_3/fa_0/a_25_6# bitslice_3/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1351 bitslice_3/fa_0/a_79_6# bitslice_3/Cin bitslice_3/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1352 bitslice_3/fa_0/a_84_6# bitslice_3/Y bitslice_3/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1353 Gnd bitslice_3/fa_0/A bitslice_3/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1354 bitslice_3/sum bitslice_3/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1355 bitslice_4/Cin bitslice_3/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1356 bitslice_3/mux21_0/nand_1/A Out3 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1357 Vdd bitslice_3/mux21_0/nand_2/B bitslice_3/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 bitslice_3/mux21_0/nand_2/a_9_6# Out3 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1359 bitslice_3/mux21_0/nand_1/A bitslice_3/mux21_0/nand_2/B bitslice_3/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1360 bitslice_3/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1361 bitslice_3/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1362 bitslice_3/fa_0/A bitslice_3/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1363 Vdd bitslice_3/mux21_0/nand_1/B bitslice_3/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 bitslice_3/mux21_0/nand_1/a_9_6# bitslice_3/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1365 bitslice_3/fa_0/A bitslice_3/mux21_0/nand_1/B bitslice_3/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1366 bitslice_3/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1367 Vdd B3 bitslice_3/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1368 bitslice_3/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1369 bitslice_3/mux21_0/nand_1/B B3 bitslice_3/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1370 Vdd A3 bitslice_3/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1371 bitslice_3/xor2_0/a_33_54# bitslice_3/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1372 bitslice_3/Y A3 bitslice_3/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1373 bitslice_3/xor2_0/a_50_54# bitslice_3/xor2_0/a_17_6# bitslice_3/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1374 Vdd subtract bitslice_3/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 bitslice_3/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1376 Gnd A3 bitslice_3/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1377 bitslice_3/xor2_0/a_33_6# bitslice_3/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1378 bitslice_3/Y bitslice_3/xor2_0/a_17_6# bitslice_3/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1379 bitslice_3/xor2_0/a_50_6# A3 bitslice_3/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1380 Gnd subtract bitslice_3/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1381 bitslice_3/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1382 Vdd inverter_0/Y bitslice_2/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1383 bitslice_2/dffpos_0/a_n19_n15# bitslice_2/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1384 bitslice_2/dffpos_0/a_n14_n84# inverter_0/Y bitslice_2/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1385 bitslice_2/dffpos_0/a_n5_n15# bitslice_2/dffpos_0/a_n34_n84# bitslice_2/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1386 Vdd bitslice_2/dffpos_0/a_n2_n86# bitslice_2/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 bitslice_2/dffpos_0/a_n2_n86# bitslice_2/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1388 bitslice_2/dffpos_0/a_25_n15# bitslice_2/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1389 bitslice_2/dffpos_0/a_30_n84# bitslice_2/dffpos_0/a_n34_n84# bitslice_2/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1390 bitslice_2/dffpos_0/a_40_n5# inverter_0/Y bitslice_2/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1391 Vdd Out2 bitslice_2/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1392 Gnd inverter_0/Y bitslice_2/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1393 Out2 bitslice_2/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1394 bitslice_2/dffpos_0/a_n19_n84# bitslice_2/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1395 bitslice_2/dffpos_0/a_n14_n84# bitslice_2/dffpos_0/a_n34_n84# bitslice_2/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1396 bitslice_2/dffpos_0/a_n5_n84# inverter_0/Y bitslice_2/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1397 Gnd bitslice_2/dffpos_0/a_n2_n86# bitslice_2/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1398 bitslice_2/dffpos_0/a_n2_n86# bitslice_2/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1399 bitslice_2/dffpos_0/a_25_n84# bitslice_2/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1400 bitslice_2/dffpos_0/a_30_n84# inverter_0/Y bitslice_2/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1401 bitslice_2/dffpos_0/a_40_n84# bitslice_2/dffpos_0/a_n34_n84# bitslice_2/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1402 Gnd Out2 bitslice_2/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 Out2 bitslice_2/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1404 Vdd bitslice_2/fa_0/A bitslice_2/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1405 bitslice_2/fa_0/a_2_74# bitslice_2/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 bitslice_2/fa_0/a_25_6# bitslice_2/Cin bitslice_2/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1407 bitslice_2/fa_0/a_33_74# bitslice_2/Y bitslice_2/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1408 Vdd bitslice_2/fa_0/A bitslice_2/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 bitslice_2/fa_0/a_46_74# bitslice_2/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1410 Vdd bitslice_2/Y bitslice_2/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 bitslice_2/fa_0/a_46_74# bitslice_2/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 bitslice_2/fa_0/a_70_6# bitslice_2/fa_0/a_25_6# bitslice_2/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1413 bitslice_2/fa_0/a_79_74# bitslice_2/Cin bitslice_2/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1414 bitslice_2/fa_0/a_84_74# bitslice_2/Y bitslice_2/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1415 Vdd bitslice_2/fa_0/A bitslice_2/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1416 bitslice_2/sum bitslice_2/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1417 bitslice_3/Cin bitslice_2/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1418 Gnd bitslice_2/fa_0/A bitslice_2/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1419 bitslice_2/fa_0/a_2_6# bitslice_2/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1420 bitslice_2/fa_0/a_25_6# bitslice_2/Cin bitslice_2/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1421 bitslice_2/fa_0/a_33_6# bitslice_2/Y bitslice_2/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1422 Gnd bitslice_2/fa_0/A bitslice_2/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 bitslice_2/fa_0/a_46_6# bitslice_2/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1424 Gnd bitslice_2/Y bitslice_2/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1425 bitslice_2/fa_0/a_46_6# bitslice_2/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1426 bitslice_2/fa_0/a_70_6# bitslice_2/fa_0/a_25_6# bitslice_2/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1427 bitslice_2/fa_0/a_79_6# bitslice_2/Cin bitslice_2/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1428 bitslice_2/fa_0/a_84_6# bitslice_2/Y bitslice_2/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1429 Gnd bitslice_2/fa_0/A bitslice_2/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 bitslice_2/sum bitslice_2/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1431 bitslice_3/Cin bitslice_2/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1432 bitslice_2/mux21_0/nand_1/A Out2 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1433 Vdd bitslice_2/mux21_0/nand_2/B bitslice_2/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1434 bitslice_2/mux21_0/nand_2/a_9_6# Out2 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1435 bitslice_2/mux21_0/nand_1/A bitslice_2/mux21_0/nand_2/B bitslice_2/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1436 bitslice_2/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1437 bitslice_2/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1438 bitslice_2/fa_0/A bitslice_2/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1439 Vdd bitslice_2/mux21_0/nand_1/B bitslice_2/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 bitslice_2/mux21_0/nand_1/a_9_6# bitslice_2/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1441 bitslice_2/fa_0/A bitslice_2/mux21_0/nand_1/B bitslice_2/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1442 bitslice_2/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1443 Vdd B2 bitslice_2/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1444 bitslice_2/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1445 bitslice_2/mux21_0/nand_1/B B2 bitslice_2/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1446 Vdd A2 bitslice_2/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1447 bitslice_2/xor2_0/a_33_54# bitslice_2/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1448 bitslice_2/Y A2 bitslice_2/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1449 bitslice_2/xor2_0/a_50_54# bitslice_2/xor2_0/a_17_6# bitslice_2/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1450 Vdd subtract bitslice_2/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1451 bitslice_2/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1452 Gnd A2 bitslice_2/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1453 bitslice_2/xor2_0/a_33_6# bitslice_2/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1454 bitslice_2/Y bitslice_2/xor2_0/a_17_6# bitslice_2/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1455 bitslice_2/xor2_0/a_50_6# A2 bitslice_2/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1456 Gnd subtract bitslice_2/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1457 bitslice_2/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1458 Vdd inverter_0/Y bitslice_1/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1459 bitslice_1/dffpos_0/a_n19_n15# bitslice_1/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1460 bitslice_1/dffpos_0/a_n14_n84# inverter_0/Y bitslice_1/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1461 bitslice_1/dffpos_0/a_n5_n15# bitslice_1/dffpos_0/a_n34_n84# bitslice_1/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1462 Vdd bitslice_1/dffpos_0/a_n2_n86# bitslice_1/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1463 bitslice_1/dffpos_0/a_n2_n86# bitslice_1/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1464 bitslice_1/dffpos_0/a_25_n15# bitslice_1/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1465 bitslice_1/dffpos_0/a_30_n84# bitslice_1/dffpos_0/a_n34_n84# bitslice_1/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1466 bitslice_1/dffpos_0/a_40_n5# inverter_0/Y bitslice_1/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1467 Vdd Out1 bitslice_1/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 Gnd inverter_0/Y bitslice_1/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1469 Out1 bitslice_1/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1470 bitslice_1/dffpos_0/a_n19_n84# bitslice_1/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1471 bitslice_1/dffpos_0/a_n14_n84# bitslice_1/dffpos_0/a_n34_n84# bitslice_1/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1472 bitslice_1/dffpos_0/a_n5_n84# inverter_0/Y bitslice_1/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1473 Gnd bitslice_1/dffpos_0/a_n2_n86# bitslice_1/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1474 bitslice_1/dffpos_0/a_n2_n86# bitslice_1/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1475 bitslice_1/dffpos_0/a_25_n84# bitslice_1/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1476 bitslice_1/dffpos_0/a_30_n84# inverter_0/Y bitslice_1/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1477 bitslice_1/dffpos_0/a_40_n84# bitslice_1/dffpos_0/a_n34_n84# bitslice_1/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1478 Gnd Out1 bitslice_1/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1479 Out1 bitslice_1/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1480 Vdd bitslice_1/fa_0/A bitslice_1/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1481 bitslice_1/fa_0/a_2_74# bitslice_1/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 bitslice_1/fa_0/a_25_6# bitslice_1/Cin bitslice_1/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1483 bitslice_1/fa_0/a_33_74# bitslice_1/Y bitslice_1/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1484 Vdd bitslice_1/fa_0/A bitslice_1/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1485 bitslice_1/fa_0/a_46_74# bitslice_1/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1486 Vdd bitslice_1/Y bitslice_1/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 bitslice_1/fa_0/a_46_74# bitslice_1/Cin Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 bitslice_1/fa_0/a_70_6# bitslice_1/fa_0/a_25_6# bitslice_1/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1489 bitslice_1/fa_0/a_79_74# bitslice_1/Cin bitslice_1/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1490 bitslice_1/fa_0/a_84_74# bitslice_1/Y bitslice_1/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1491 Vdd bitslice_1/fa_0/A bitslice_1/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1492 bitslice_1/sum bitslice_1/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1493 bitslice_2/Cin bitslice_1/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1494 Gnd bitslice_1/fa_0/A bitslice_1/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1495 bitslice_1/fa_0/a_2_6# bitslice_1/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 bitslice_1/fa_0/a_25_6# bitslice_1/Cin bitslice_1/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1497 bitslice_1/fa_0/a_33_6# bitslice_1/Y bitslice_1/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1498 Gnd bitslice_1/fa_0/A bitslice_1/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1499 bitslice_1/fa_0/a_46_6# bitslice_1/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1500 Gnd bitslice_1/Y bitslice_1/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 bitslice_1/fa_0/a_46_6# bitslice_1/Cin Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1502 bitslice_1/fa_0/a_70_6# bitslice_1/fa_0/a_25_6# bitslice_1/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1503 bitslice_1/fa_0/a_79_6# bitslice_1/Cin bitslice_1/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1504 bitslice_1/fa_0/a_84_6# bitslice_1/Y bitslice_1/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1505 Gnd bitslice_1/fa_0/A bitslice_1/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 bitslice_1/sum bitslice_1/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1507 bitslice_2/Cin bitslice_1/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1508 bitslice_1/mux21_0/nand_1/A Out1 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1509 Vdd bitslice_1/mux21_0/nand_2/B bitslice_1/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 bitslice_1/mux21_0/nand_2/a_9_6# Out1 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1511 bitslice_1/mux21_0/nand_1/A bitslice_1/mux21_0/nand_2/B bitslice_1/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1512 bitslice_1/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1513 bitslice_1/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1514 bitslice_1/fa_0/A bitslice_1/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1515 Vdd bitslice_1/mux21_0/nand_1/B bitslice_1/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 bitslice_1/mux21_0/nand_1/a_9_6# bitslice_1/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1517 bitslice_1/fa_0/A bitslice_1/mux21_0/nand_1/B bitslice_1/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1518 bitslice_1/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1519 Vdd B1 bitslice_1/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1520 bitslice_1/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1521 bitslice_1/mux21_0/nand_1/B B1 bitslice_1/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1522 Vdd A1 bitslice_1/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1523 bitslice_1/xor2_0/a_33_54# bitslice_1/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1524 bitslice_1/Y A1 bitslice_1/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1525 bitslice_1/xor2_0/a_50_54# bitslice_1/xor2_0/a_17_6# bitslice_1/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1526 Vdd subtract bitslice_1/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1527 bitslice_1/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1528 Gnd A1 bitslice_1/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1529 bitslice_1/xor2_0/a_33_6# bitslice_1/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1530 bitslice_1/Y bitslice_1/xor2_0/a_17_6# bitslice_1/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1531 bitslice_1/xor2_0/a_50_6# A1 bitslice_1/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1532 Gnd subtract bitslice_1/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1533 bitslice_1/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1534 Vdd inverter_0/Y bitslice_0/dffpos_0/a_n34_n84# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1535 bitslice_0/dffpos_0/a_n19_n15# bitslice_0/sum Vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1536 bitslice_0/dffpos_0/a_n14_n84# inverter_0/Y bitslice_0/dffpos_0/a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1537 bitslice_0/dffpos_0/a_n5_n15# bitslice_0/dffpos_0/a_n34_n84# bitslice_0/dffpos_0/a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1538 Vdd bitslice_0/dffpos_0/a_n2_n86# bitslice_0/dffpos_0/a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1539 bitslice_0/dffpos_0/a_n2_n86# bitslice_0/dffpos_0/a_n14_n84# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1540 bitslice_0/dffpos_0/a_25_n15# bitslice_0/dffpos_0/a_n2_n86# Vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1541 bitslice_0/dffpos_0/a_30_n84# bitslice_0/dffpos_0/a_n34_n84# bitslice_0/dffpos_0/a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1542 bitslice_0/dffpos_0/a_40_n5# inverter_0/Y bitslice_0/dffpos_0/a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1543 Vdd Out0 bitslice_0/dffpos_0/a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1544 Gnd inverter_0/Y bitslice_0/dffpos_0/a_n34_n84# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1545 Out0 bitslice_0/dffpos_0/a_30_n84# Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1546 bitslice_0/dffpos_0/a_n19_n84# bitslice_0/sum Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1547 bitslice_0/dffpos_0/a_n14_n84# bitslice_0/dffpos_0/a_n34_n84# bitslice_0/dffpos_0/a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1548 bitslice_0/dffpos_0/a_n5_n84# inverter_0/Y bitslice_0/dffpos_0/a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1549 Gnd bitslice_0/dffpos_0/a_n2_n86# bitslice_0/dffpos_0/a_n5_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1550 bitslice_0/dffpos_0/a_n2_n86# bitslice_0/dffpos_0/a_n14_n84# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1551 bitslice_0/dffpos_0/a_25_n84# bitslice_0/dffpos_0/a_n2_n86# Gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1552 bitslice_0/dffpos_0/a_30_n84# inverter_0/Y bitslice_0/dffpos_0/a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1553 bitslice_0/dffpos_0/a_40_n84# bitslice_0/dffpos_0/a_n34_n84# bitslice_0/dffpos_0/a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1554 Gnd Out0 bitslice_0/dffpos_0/a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1555 Out0 bitslice_0/dffpos_0/a_30_n84# Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1556 Vdd bitslice_0/fa_0/A bitslice_0/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1557 bitslice_0/fa_0/a_2_74# bitslice_0/Y Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1558 bitslice_0/fa_0/a_25_6# subtract bitslice_0/fa_0/a_2_74# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1559 bitslice_0/fa_0/a_33_74# bitslice_0/Y bitslice_0/fa_0/a_25_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1560 Vdd bitslice_0/fa_0/A bitslice_0/fa_0/a_33_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1561 bitslice_0/fa_0/a_46_74# bitslice_0/fa_0/A Vdd Vdd pfet w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1562 Vdd bitslice_0/Y bitslice_0/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 bitslice_0/fa_0/a_46_74# subtract Vdd Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1564 bitslice_0/fa_0/a_70_6# bitslice_0/fa_0/a_25_6# bitslice_0/fa_0/a_46_74# Vdd pfet w=20 l=2
+  ad=140 pd=54 as=0 ps=0
M1565 bitslice_0/fa_0/a_79_74# subtract bitslice_0/fa_0/a_70_6# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1566 bitslice_0/fa_0/a_84_74# bitslice_0/Y bitslice_0/fa_0/a_79_74# Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1567 Vdd bitslice_0/fa_0/A bitslice_0/fa_0/a_84_74# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1568 bitslice_0/sum bitslice_0/fa_0/a_70_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1569 bitslice_1/Cin bitslice_0/fa_0/a_25_6# Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1570 Gnd bitslice_0/fa_0/A bitslice_0/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=110 ps=62
M1571 bitslice_0/fa_0/a_2_6# bitslice_0/Y Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1572 bitslice_0/fa_0/a_25_6# subtract bitslice_0/fa_0/a_2_6# Gnd nfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1573 bitslice_0/fa_0/a_33_6# bitslice_0/Y bitslice_0/fa_0/a_25_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1574 Gnd bitslice_0/fa_0/A bitslice_0/fa_0/a_33_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1575 bitslice_0/fa_0/a_46_6# bitslice_0/fa_0/A Gnd Gnd nfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1576 Gnd bitslice_0/Y bitslice_0/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 bitslice_0/fa_0/a_46_6# subtract Gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1578 bitslice_0/fa_0/a_70_6# bitslice_0/fa_0/a_25_6# bitslice_0/fa_0/a_46_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1579 bitslice_0/fa_0/a_79_6# subtract bitslice_0/fa_0/a_70_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1580 bitslice_0/fa_0/a_84_6# bitslice_0/Y bitslice_0/fa_0/a_79_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1581 Gnd bitslice_0/fa_0/A bitslice_0/fa_0/a_84_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1582 bitslice_0/sum bitslice_0/fa_0/a_70_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1583 bitslice_1/Cin bitslice_0/fa_0/a_25_6# Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1584 bitslice_0/mux21_0/nand_1/A Out0 Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1585 Vdd bitslice_0/mux21_0/nand_2/B bitslice_0/mux21_0/nand_1/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1586 bitslice_0/mux21_0/nand_2/a_9_6# Out0 Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1587 bitslice_0/mux21_0/nand_1/A bitslice_0/mux21_0/nand_2/B bitslice_0/mux21_0/nand_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1588 bitslice_0/mux21_0/nand_2/B loadB Vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1589 bitslice_0/mux21_0/nand_2/B loadB Gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1590 bitslice_0/fa_0/A bitslice_0/mux21_0/nand_1/A Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1591 Vdd bitslice_0/mux21_0/nand_1/B bitslice_0/fa_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 bitslice_0/mux21_0/nand_1/a_9_6# bitslice_0/mux21_0/nand_1/A Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1593 bitslice_0/fa_0/A bitslice_0/mux21_0/nand_1/B bitslice_0/mux21_0/nand_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1594 bitslice_0/mux21_0/nand_1/B loadB Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1595 Vdd B0 bitslice_0/mux21_0/nand_1/B Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1596 bitslice_0/mux21_0/nand_0/a_9_6# loadB Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1597 bitslice_0/mux21_0/nand_1/B B0 bitslice_0/mux21_0/nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1598 Vdd A0 bitslice_0/xor2_0/a_17_6# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1599 bitslice_0/xor2_0/a_33_54# bitslice_0/xor2_0/a_28_44# Vdd Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1600 bitslice_0/Y A0 bitslice_0/xor2_0/a_33_54# Vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1601 bitslice_0/xor2_0/a_50_54# bitslice_0/xor2_0/a_17_6# bitslice_0/Y Vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1602 Vdd subtract bitslice_0/xor2_0/a_50_54# Vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1603 bitslice_0/xor2_0/a_28_44# subtract Vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1604 Gnd A0 bitslice_0/xor2_0/a_17_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100 ps=50
M1605 bitslice_0/xor2_0/a_33_6# bitslice_0/xor2_0/a_28_44# Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1606 bitslice_0/Y bitslice_0/xor2_0/a_17_6# bitslice_0/xor2_0/a_33_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1607 bitslice_0/xor2_0/a_50_6# A0 bitslice_0/Y Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1608 Gnd subtract bitslice_0/xor2_0/a_50_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1609 bitslice_0/xor2_0/a_28_44# subtract Gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1610 inverter_0/A loadR Vdd Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1611 Vdd clk inverter_0/A Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1612 nand_0/a_9_6# loadR Gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1613 inverter_0/A clk nand_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 bitslice_2/fa_0/a_70_6# bitslice_2/Cin 2.233260fF
C1 bitslice_3/mux21_0/nand_2/B Vdd 5.855850fF
C2 bitslice_1/mux21_0/nand_1/B Vdd 2.097720fF
C3 Vdd bitslice_1/xor2_0/a_17_6# 2.059560fF
C4 bitslice_4/dffpos_0/a_n34_n84# bitslice_4/dffpos_0/a_30_n84# 2.081040fF
C5 bitslice_3/dffpos_0/a_n34_n84# inverter_0/Y 2.571480fF
C6 inverter_0/Y bitslice_3/dffpos_0/a_n2_n86# 3.159600fF
C7 bitslice_5/dffpos_0/a_30_n84# bitslice_5/dffpos_0/a_n34_n84# 2.081040fF
C8 bitslice_7/Cin bitslice_7/fa_0/a_70_6# 2.233260fF
C9 Vdd bitslice_5/fa_0/A 8.476560fF
C10 bitslice_1/sum Gnd 5.857320fF
C11 loadB subtract 2.514300fF
C12 inverter_0/Y bitslice_0/dffpos_0/a_n34_n84# 2.571480fF
C13 bitslice_1/xor2_0/a_28_44# Vdd 2.119800fF
C14 Vdd bitslice_3/fa_0/A 8.476560fF
C15 inverter_0/Y bitslice_0/dffpos_0/a_n2_n86# 3.159600fF
C16 inverter_0/Y Gnd 2.544000fF
C17 loadB Gnd 5.499840fF
C18 bitslice_4/mux21_0/nand_1/B Vdd 2.097720fF
C19 bitslice_6/dffpos_0/a_30_n84# bitslice_6/dffpos_0/a_n34_n84# 2.081040fF
C20 bitslice_4/fa_0/a_70_6# bitslice_4/Cin 2.233260fF
C21 Gnd bitslice_0/sum 5.857320fF
C22 bitslice_3/fa_0/a_70_6# bitslice_3/Cin 2.233260fF
C23 bitslice_4/dffpos_0/a_n2_n86# inverter_0/Y 3.159600fF
C24 bitslice_6/sum Gnd 5.857320fF
C25 subtract bitslice_0/fa_0/a_70_6# 2.233260fF
C26 bitslice_5/fa_0/a_25_6# Vdd 3.134880fF
C27 bitslice_2/sum Gnd 5.857320fF
C28 Vdd bitslice_7/xor2_0/a_17_6# 2.059560fF
C29 bitslice_6/mux21_0/nand_2/B Vdd 5.855850fF
C30 inverter_0/Y bitslice_7/dffpos_0/a_n34_n84# 2.571480fF
C31 bitslice_7/dffpos_0/a_n34_n84# bitslice_7/dffpos_0/a_30_n84# 2.081040fF
C32 bitslice_0/dffpos_0/a_30_n84# bitslice_0/dffpos_0/a_n34_n84# 2.081040fF
C33 Vdd bitslice_2/fa_0/a_25_6# 3.134880fF
C34 Vdd bitslice_0/xor2_0/a_17_6# 2.059560fF
C35 inverter_0/Y bitslice_2/dffpos_0/a_n2_n86# 3.159600fF
C36 Vdd bitslice_0/xor2_0/a_28_44# 2.119800fF
C37 Vdd bitslice_2/fa_0/A 8.476560fF
C38 bitslice_2/mux21_0/nand_2/B Vdd 5.855850fF
C39 bitslice_6/fa_0/A Vdd 8.476560fF
C40 Gnd subtract 3.855720fF
C41 bitslice_2/dffpos_0/a_30_n84# bitslice_2/dffpos_0/a_n34_n84# 2.081040fF
C42 Vdd bitslice_3/xor2_0/a_28_44# 2.119800fF
C43 bitslice_7/xor2_0/a_28_44# Vdd 2.119800fF
C44 bitslice_3/dffpos_0/a_30_n84# bitslice_3/dffpos_0/a_n34_n84# 2.081040fF
C45 inverter_0/Y bitslice_5/dffpos_0/a_n34_n84# 2.571480fF
C46 inverter_0/Y bitslice_1/dffpos_0/a_n2_n86# 3.159600fF
C47 inverter_0/Y bitslice_5/dffpos_0/a_n2_n86# 3.159600fF
C48 Gnd bitslice_3/sum 5.857320fF
C49 bitslice_5/xor2_0/a_28_44# Vdd 2.119800fF
C50 bitslice_3/fa_0/a_25_6# Vdd 3.134880fF
C51 Gnd bitslice_4/sum 5.857320fF
C52 bitslice_5/xor2_0/a_17_6# Vdd 2.059560fF
C53 inverter_0/Y Vdd 11.673119fF
C54 inverter_0/Y bitslice_2/dffpos_0/a_n34_n84# 2.571480fF
C55 bitslice_5/mux21_0/nand_2/B Vdd 5.855850fF
C56 inverter_0/Y bitslice_7/dffpos_0/a_n2_n86# 3.159600fF
C57 loadB Vdd 6.672270fF
C58 bitslice_7/fa_0/A Vdd 8.476560fF
C59 bitslice_1/mux21_0/nand_2/B Vdd 5.855850fF
C60 inverter_0/Y bitslice_6/dffpos_0/a_n2_n86# 3.159600fF
C61 bitslice_6/xor2_0/a_28_44# Vdd 2.119800fF
C62 bitslice_4/fa_0/a_25_6# Vdd 3.134880fF
C63 inverter_0/Y bitslice_6/dffpos_0/a_n34_n84# 2.571480fF
C64 bitslice_7/mux21_0/nand_2/B Vdd 5.855850fF
C65 bitslice_6/mux21_0/nand_1/B Vdd 2.097720fF
C66 Vdd bitslice_0/fa_0/a_25_6# 3.134880fF
C67 bitslice_1/fa_0/A Vdd 8.476560fF
C68 bitslice_5/sum Gnd 5.857320fF
C69 Vdd bitslice_3/xor2_0/a_17_6# 2.059560fF
C70 bitslice_7/fa_0/a_25_6# Vdd 3.134880fF
C71 bitslice_1/dffpos_0/a_30_n84# bitslice_1/dffpos_0/a_n34_n84# 2.081040fF
C72 Vdd bitslice_0/mux21_0/nand_2/B 5.855850fF
C73 bitslice_4/fa_0/A Vdd 8.476560fF
C74 bitslice_2/xor2_0/a_17_6# Vdd 2.059560fF
C75 bitslice_1/Cin bitslice_1/fa_0/a_70_6# 2.233260fF
C76 subtract Vdd 6.123960fF
C77 Vdd bitslice_7/mux21_0/nand_1/B 2.097720fF
C78 bitslice_6/fa_0/a_25_6# Vdd 3.134880fF
C79 gundy Gnd 5.857320fF
C80 bitslice_6/xor2_0/a_17_6# Vdd 2.059560fF
C81 Vdd bitslice_3/mux21_0/nand_1/B 2.097720fF
C82 bitslice_5/mux21_0/nand_1/B Vdd 2.097720fF
C83 Vdd bitslice_2/xor2_0/a_28_44# 2.119800fF
C84 Gnd Vdd 4.961880fF
C85 bitslice_4/dffpos_0/a_n34_n84# inverter_0/Y 2.571480fF
C86 Vdd bitslice_1/fa_0/a_25_6# 3.134880fF
C87 bitslice_4/xor2_0/a_28_44# Vdd 2.119800fF
C88 bitslice_4/mux21_0/nand_2/B Vdd 5.855850fF
C89 bitslice_6/fa_0/a_70_6# bitslice_6/Cin 2.233260fF
C90 Vdd bitslice_0/fa_0/A 8.476560fF
C91 bitslice_2/mux21_0/nand_1/B Vdd 2.097720fF
C92 bitslice_4/xor2_0/a_17_6# Vdd 2.059560fF
C93 Vdd bitslice_0/mux21_0/nand_1/B 2.097720fF
C94 inverter_0/Y bitslice_1/dffpos_0/a_n34_n84# 2.571480fF
C95 bitslice_5/fa_0/a_70_6# bitslice_5/Cin 2.233260fF
C96 bitslice_0/Y gnd! 18.021119fF
C97 bitslice_0/xor2_0/a_17_6# gnd! 4.666380fF
C98 bitslice_0/xor2_0/a_28_44# gnd! 4.104630fF
C99 bitslice_0/fa_0/A gnd! 7.718120fF
C100 bitslice_0/mux21_0/nand_1/B gnd! 3.001320fF
C101 bitslice_0/mux21_0/nand_1/A gnd! 6.037200fF
C102 bitslice_0/mux21_0/nand_2/B gnd! 2.145240fF
C103 Out0 gnd! 87.604953fF
C104 bitslice_0/sum gnd! 8.877960fF
C105 bitslice_0/fa_0/a_70_6# gnd! 3.242790fF
C106 bitslice_0/fa_0/a_25_6# gnd! 9.314280fF
C107 bitslice_0/dffpos_0/a_30_n84# gnd! 3.784590fF
C108 bitslice_0/dffpos_0/a_n14_n84# gnd! 4.801770fF
C109 bitslice_0/dffpos_0/a_n2_n86# gnd! 5.164560fF
C110 bitslice_0/dffpos_0/a_n34_n84# gnd! 8.655120fF
C111 bitslice_1/Y gnd! 18.021119fF
C112 bitslice_1/xor2_0/a_17_6# gnd! 4.666380fF
C113 bitslice_1/xor2_0/a_28_44# gnd! 4.104630fF
C114 bitslice_1/fa_0/A gnd! 7.718120fF
C115 bitslice_1/mux21_0/nand_1/B gnd! 3.001320fF
C116 bitslice_1/mux21_0/nand_1/A gnd! 6.037200fF
C117 bitslice_1/mux21_0/nand_2/B gnd! 2.145240fF
C118 Out1 gnd! 76.024156fF
C119 bitslice_1/sum gnd! 8.877960fF
C120 bitslice_1/fa_0/a_70_6# gnd! 3.242790fF
C121 bitslice_1/fa_0/a_25_6# gnd! 9.314280fF
C122 bitslice_1/dffpos_0/a_30_n84# gnd! 3.784590fF
C123 bitslice_1/dffpos_0/a_n14_n84# gnd! 4.801770fF
C124 bitslice_1/dffpos_0/a_n2_n86# gnd! 5.164560fF
C125 bitslice_1/dffpos_0/a_n34_n84# gnd! 8.655120fF
C126 bitslice_2/Y gnd! 18.021119fF
C127 bitslice_2/xor2_0/a_17_6# gnd! 4.666380fF
C128 bitslice_2/xor2_0/a_28_44# gnd! 4.104630fF
C129 bitslice_2/fa_0/A gnd! 7.718120fF
C130 bitslice_2/mux21_0/nand_1/B gnd! 3.001320fF
C131 bitslice_2/mux21_0/nand_1/A gnd! 6.037200fF
C132 bitslice_2/mux21_0/nand_2/B gnd! 2.145240fF
C133 Out2 gnd! 67.891609fF
C134 bitslice_2/sum gnd! 8.877960fF
C135 bitslice_2/fa_0/a_70_6# gnd! 3.242790fF
C136 bitslice_2/fa_0/a_25_6# gnd! 9.314280fF
C137 bitslice_2/dffpos_0/a_30_n84# gnd! 3.784590fF
C138 bitslice_2/dffpos_0/a_n14_n84# gnd! 4.801770fF
C139 bitslice_2/dffpos_0/a_n2_n86# gnd! 5.164560fF
C140 bitslice_2/dffpos_0/a_n34_n84# gnd! 8.655120fF
C141 bitslice_3/Y gnd! 18.021119fF
C142 bitslice_3/xor2_0/a_17_6# gnd! 4.666380fF
C143 bitslice_3/xor2_0/a_28_44# gnd! 4.104630fF
C144 bitslice_3/fa_0/A gnd! 7.718120fF
C145 bitslice_3/mux21_0/nand_1/B gnd! 3.001320fF
C146 bitslice_3/mux21_0/nand_1/A gnd! 6.037200fF
C147 bitslice_3/mux21_0/nand_2/B gnd! 2.145240fF
C148 Out3 gnd! 58.928160fF
C149 bitslice_3/sum gnd! 8.877960fF
C150 bitslice_3/fa_0/a_70_6# gnd! 3.242790fF
C151 bitslice_3/fa_0/a_25_6# gnd! 9.314280fF
C152 bitslice_3/dffpos_0/a_30_n84# gnd! 3.784590fF
C153 bitslice_3/dffpos_0/a_n14_n84# gnd! 4.801770fF
C154 bitslice_3/dffpos_0/a_n2_n86# gnd! 5.164560fF
C155 bitslice_3/dffpos_0/a_n34_n84# gnd! 8.655120fF
C156 bitslice_4/Y gnd! 18.021119fF
C157 bitslice_4/xor2_0/a_17_6# gnd! 4.666380fF
C158 bitslice_4/xor2_0/a_28_44# gnd! 4.104630fF
C159 bitslice_4/fa_0/A gnd! 7.718120fF
C160 bitslice_4/mux21_0/nand_1/B gnd! 3.001320fF
C161 bitslice_4/mux21_0/nand_1/A gnd! 6.037200fF
C162 bitslice_4/mux21_0/nand_2/B gnd! 2.145240fF
C163 Out4 gnd! 50.394660fF
C164 bitslice_4/sum gnd! 8.877960fF
C165 bitslice_4/fa_0/a_70_6# gnd! 3.242790fF
C166 bitslice_4/fa_0/a_25_6# gnd! 9.314280fF
C167 bitslice_4/dffpos_0/a_30_n84# gnd! 3.784590fF
C168 bitslice_4/dffpos_0/a_n14_n84# gnd! 4.801770fF
C169 bitslice_4/dffpos_0/a_n2_n86# gnd! 5.164560fF
C170 bitslice_4/dffpos_0/a_n34_n84# gnd! 8.655120fF
C171 bitslice_5/Y gnd! 18.021119fF
C172 bitslice_5/xor2_0/a_17_6# gnd! 4.666380fF
C173 bitslice_5/xor2_0/a_28_44# gnd! 4.104630fF
C174 bitslice_5/fa_0/A gnd! 7.718120fF
C175 bitslice_5/mux21_0/nand_1/B gnd! 3.001320fF
C176 bitslice_5/mux21_0/nand_1/A gnd! 6.037200fF
C177 bitslice_5/mux21_0/nand_2/B gnd! 2.145240fF
C178 Out5 gnd! 41.783863fF
C179 bitslice_5/sum gnd! 8.877960fF
C180 bitslice_5/fa_0/a_70_6# gnd! 3.242790fF
C181 bitslice_5/fa_0/a_25_6# gnd! 9.314280fF
C182 bitslice_5/dffpos_0/a_30_n84# gnd! 3.784590fF
C183 bitslice_5/dffpos_0/a_n14_n84# gnd! 4.801770fF
C184 bitslice_5/dffpos_0/a_n2_n86# gnd! 5.164560fF
C185 bitslice_5/dffpos_0/a_n34_n84# gnd! 8.655120fF
C186 bitslice_6/Y gnd! 18.021119fF
C187 bitslice_6/xor2_0/a_17_6# gnd! 4.666380fF
C188 bitslice_6/xor2_0/a_28_44# gnd! 4.104630fF
C189 bitslice_6/fa_0/A gnd! 7.718120fF
C190 bitslice_6/mux21_0/nand_1/B gnd! 3.001320fF
C191 bitslice_6/mux21_0/nand_1/A gnd! 6.037200fF
C192 bitslice_6/mux21_0/nand_2/B gnd! 2.145240fF
C193 Out6 gnd! 33.352602fF
C194 bitslice_6/sum gnd! 8.877960fF
C195 bitslice_6/fa_0/a_70_6# gnd! 3.242790fF
C196 bitslice_6/fa_0/a_25_6# gnd! 9.314280fF
C197 bitslice_6/dffpos_0/a_30_n84# gnd! 3.784590fF
C198 bitslice_6/dffpos_0/a_n14_n84# gnd! 4.801770fF
C199 bitslice_6/dffpos_0/a_n2_n86# gnd! 5.164560fF
C200 bitslice_6/dffpos_0/a_n34_n84# gnd! 8.655120fF
C201 Gnd gnd! 1242.410750fF
C202 bitslice_7/Y gnd! 18.021119fF
C203 subtract gnd! 101.129359fF
C204 bitslice_7/xor2_0/a_17_6# gnd! 4.666380fF
C205 bitslice_7/xor2_0/a_28_44# gnd! 4.104630fF
C206 loadB gnd! 155.956141fF
C207 bitslice_7/fa_0/A gnd! 7.718120fF
C208 bitslice_7/mux21_0/nand_1/B gnd! 3.001320fF
C209 bitslice_7/mux21_0/nand_1/A gnd! 6.037200fF
C210 bitslice_7/mux21_0/nand_2/B gnd! 2.145240fF
C211 Out7 gnd! 25.139992fF
C212 bitslice_7/fa_0/a_70_6# gnd! 3.242790fF
C213 bitslice_7/fa_0/a_25_6# gnd! 9.314280fF
C214 bitslice_7/dffpos_0/a_30_n84# gnd! 3.784590fF
C215 bitslice_7/dffpos_0/a_n14_n84# gnd! 4.801770fF
C216 bitslice_7/dffpos_0/a_n2_n86# gnd! 5.164560fF
C217 bitslice_7/dffpos_0/a_n34_n84# gnd! 8.655120fF
C218 inverter_0/Y gnd! 148.452219fF
C219 inverter_0/A gnd! 8.251561fF
