* SPICE3 file created from dffpos.ext - technology: scmos

.option scale=0.3u

M1000 vdd a_n33_n56# clk Vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1001 a_n19_n15# D vdd Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1002 a_n14_n84# a_n33_n56# a_n19_n15# Vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1003 a_n5_n15# clk a_n14_n84# Vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1004 vdd a_n2_n86# a_n5_n15# Vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_n2_n86# a_n14_n84# vdd Vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 a_25_n15# a_n2_n86# vdd Vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1007 a_30_n84# clk a_25_n15# Vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1008 a_40_n5# a_n33_n56# a_30_n84# Vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1009 vdd Q a_40_n5# Vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_n27_n84# a_n33_n56# clk Gnd nfet w=20 l=2
+  ad=110 pd=52 as=100 ps=50
M1011 Q a_30_n84# vdd Vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1012 a_n19_n84# D a_n27_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1013 a_n14_n84# clk a_n19_n84# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1014 a_n5_n84# a_n33_n56# a_n14_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1015 gnd a_n2_n86# a_n5_n84# Gnd nfet w=10 l=2
+  ad=230 pd=116 as=0 ps=0
M1016 a_n2_n86# a_n14_n84# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1017 a_25_n84# a_n2_n86# gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1018 a_30_n84# a_n33_n56# a_25_n84# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1019 a_40_n84# clk a_30_n84# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1020 gnd Q a_40_n84# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 Q a_30_n84# gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 a_30_n84# clk 2.081040fF
C1 a_n33_n56# a_n2_n86# 3.159600fF
C2 a_n33_n56# clk 2.571480fF
C3 gnd gnd! 7.687800fF
C4 a_30_n84# gnd! 3.784590fF
C5 Q gnd! 6.264360fF
C6 a_n14_n84# gnd! 5.061090fF
C7 a_n2_n86# gnd! 5.385720fF
C8 clk gnd! 9.404880fF
C9 a_n33_n56# gnd! 12.488580fF
C10 vdd gnd! 9.030600fF
