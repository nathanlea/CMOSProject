* FILE: mux21.sp

********************** begin header *****************************

* Sample Spice Header file for Generic 2.5V 0.25 um process (mmi25)

.OPTIONS post NOMOD post_version=9601

**################################################
* Only Typical/Typical spice models included
.include '${MMI_TOOLS}/sue/schematics/mspice/mmi25.mod'
* NOTE: these are contrived spice models
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=0,2,10,12 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3,13 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.6u
.param lp_min   =  0.6u

* used in source/drain area/perimeter calculation
.param sdd        =  0.66

.PARAM vddp=2.25	$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 5p 10n

*********************** end header ******************************

* SPICE netlist for "mux21" generated by MMI_SUE5.6.18 on Sun Nov 08 
*+ 19:30:07 CST 2015.

* start main CELL mux21
* .SUBCKT mux21 In_0 In_1 Out Sel Sel_bar 
M_1 Out Sel In_1 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_2 Out Sel_bar In_1 vdd p W='3*1u' L=lp_min ad='areap(3,sdd)' 
+ as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
M_3 Out Sel_bar In_0 gnd n W='3*1u' L=ln_min ad='arean(3,sdd)' 
+ as='arean(3,sdd)' pd='perin(3,sdd)' ps='perin(3,sdd)' 
M_4 Out Sel In_0 vdd p W='3*1u' L=lp_min ad='areap(3,sdd)' 
+ as='areap(3,sdd)' pd='perip(3,sdd)' ps='perip(3,sdd)' 
* .ENDS	$ mux21

.END

